module laplacian (CLK,
    rst,
    valid_in,
    valid_out,
    pixel_in,
    pixel_out);
 input CLK;
 input rst;
 input valid_in;
 output valid_out;
 input [7:0] pixel_in;
 output [7:0] pixel_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire \col_input[0] ;
 wire \col_input[10] ;
 wire \col_input[11] ;
 wire \col_input[12] ;
 wire \col_input[13] ;
 wire \col_input[14] ;
 wire \col_input[15] ;
 wire \col_input[16] ;
 wire \col_input[17] ;
 wire \col_input[18] ;
 wire \col_input[19] ;
 wire \col_input[1] ;
 wire \col_input[20] ;
 wire \col_input[21] ;
 wire \col_input[22] ;
 wire \col_input[23] ;
 wire \col_input[24] ;
 wire \col_input[25] ;
 wire \col_input[26] ;
 wire \col_input[27] ;
 wire \col_input[28] ;
 wire \col_input[29] ;
 wire \col_input[2] ;
 wire \col_input[30] ;
 wire \col_input[31] ;
 wire \col_input[3] ;
 wire \col_input[4] ;
 wire \col_input[5] ;
 wire \col_input[6] ;
 wire \col_input[7] ;
 wire \col_input[8] ;
 wire \col_input[9] ;
 wire \col_operation[0] ;
 wire \col_operation[1] ;
 wire \col_operation[2] ;
 wire \col_operation[3] ;
 wire \col_operation[4] ;
 wire \first_row[0][0] ;
 wire \first_row[0][1] ;
 wire \first_row[0][2] ;
 wire \first_row[0][3] ;
 wire \first_row[0][4] ;
 wire \first_row[0][5] ;
 wire \first_row[0][6] ;
 wire \first_row[0][7] ;
 wire \first_row[10][0] ;
 wire \first_row[10][1] ;
 wire \first_row[10][2] ;
 wire \first_row[10][3] ;
 wire \first_row[10][4] ;
 wire \first_row[10][5] ;
 wire \first_row[10][6] ;
 wire \first_row[10][7] ;
 wire \first_row[11][0] ;
 wire \first_row[11][1] ;
 wire \first_row[11][2] ;
 wire \first_row[11][3] ;
 wire \first_row[11][4] ;
 wire \first_row[11][5] ;
 wire \first_row[11][6] ;
 wire \first_row[11][7] ;
 wire \first_row[12][0] ;
 wire \first_row[12][1] ;
 wire \first_row[12][2] ;
 wire \first_row[12][3] ;
 wire \first_row[12][4] ;
 wire \first_row[12][5] ;
 wire \first_row[12][6] ;
 wire \first_row[12][7] ;
 wire \first_row[13][0] ;
 wire \first_row[13][1] ;
 wire \first_row[13][2] ;
 wire \first_row[13][3] ;
 wire \first_row[13][4] ;
 wire \first_row[13][5] ;
 wire \first_row[13][6] ;
 wire \first_row[13][7] ;
 wire \first_row[14][0] ;
 wire \first_row[14][1] ;
 wire \first_row[14][2] ;
 wire \first_row[14][3] ;
 wire \first_row[14][4] ;
 wire \first_row[14][5] ;
 wire \first_row[14][6] ;
 wire \first_row[14][7] ;
 wire \first_row[15][0] ;
 wire \first_row[15][1] ;
 wire \first_row[15][2] ;
 wire \first_row[15][3] ;
 wire \first_row[15][4] ;
 wire \first_row[15][5] ;
 wire \first_row[15][6] ;
 wire \first_row[15][7] ;
 wire \first_row[16][0] ;
 wire \first_row[16][1] ;
 wire \first_row[16][2] ;
 wire \first_row[16][3] ;
 wire \first_row[16][4] ;
 wire \first_row[16][5] ;
 wire \first_row[16][6] ;
 wire \first_row[16][7] ;
 wire \first_row[17][0] ;
 wire \first_row[17][1] ;
 wire \first_row[17][2] ;
 wire \first_row[17][3] ;
 wire \first_row[17][4] ;
 wire \first_row[17][5] ;
 wire \first_row[17][6] ;
 wire \first_row[17][7] ;
 wire \first_row[1][0] ;
 wire \first_row[1][1] ;
 wire \first_row[1][2] ;
 wire \first_row[1][3] ;
 wire \first_row[1][4] ;
 wire \first_row[1][5] ;
 wire \first_row[1][6] ;
 wire \first_row[1][7] ;
 wire \first_row[2][0] ;
 wire \first_row[2][1] ;
 wire \first_row[2][2] ;
 wire \first_row[2][3] ;
 wire \first_row[2][4] ;
 wire \first_row[2][5] ;
 wire \first_row[2][6] ;
 wire \first_row[2][7] ;
 wire \first_row[3][0] ;
 wire \first_row[3][1] ;
 wire \first_row[3][2] ;
 wire \first_row[3][3] ;
 wire \first_row[3][4] ;
 wire \first_row[3][5] ;
 wire \first_row[3][6] ;
 wire \first_row[3][7] ;
 wire \first_row[4][0] ;
 wire \first_row[4][1] ;
 wire \first_row[4][2] ;
 wire \first_row[4][3] ;
 wire \first_row[4][4] ;
 wire \first_row[4][5] ;
 wire \first_row[4][6] ;
 wire \first_row[4][7] ;
 wire \first_row[5][0] ;
 wire \first_row[5][1] ;
 wire \first_row[5][2] ;
 wire \first_row[5][3] ;
 wire \first_row[5][4] ;
 wire \first_row[5][5] ;
 wire \first_row[5][6] ;
 wire \first_row[5][7] ;
 wire \first_row[6][0] ;
 wire \first_row[6][1] ;
 wire \first_row[6][2] ;
 wire \first_row[6][3] ;
 wire \first_row[6][4] ;
 wire \first_row[6][5] ;
 wire \first_row[6][6] ;
 wire \first_row[6][7] ;
 wire \first_row[7][0] ;
 wire \first_row[7][1] ;
 wire \first_row[7][2] ;
 wire \first_row[7][3] ;
 wire \first_row[7][4] ;
 wire \first_row[7][5] ;
 wire \first_row[7][6] ;
 wire \first_row[7][7] ;
 wire \first_row[8][0] ;
 wire \first_row[8][1] ;
 wire \first_row[8][2] ;
 wire \first_row[8][3] ;
 wire \first_row[8][4] ;
 wire \first_row[8][5] ;
 wire \first_row[8][6] ;
 wire \first_row[8][7] ;
 wire \first_row[9][0] ;
 wire \first_row[9][1] ;
 wire \first_row[9][2] ;
 wire \first_row[9][3] ;
 wire \first_row[9][4] ;
 wire \first_row[9][5] ;
 wire \first_row[9][6] ;
 wire \first_row[9][7] ;
 wire \k[0] ;
 wire \k[10] ;
 wire \k[11] ;
 wire \k[12] ;
 wire \k[13] ;
 wire \k[14] ;
 wire \k[15] ;
 wire \k[16] ;
 wire \k[17] ;
 wire \k[18] ;
 wire \k[19] ;
 wire \k[1] ;
 wire \k[20] ;
 wire \k[21] ;
 wire \k[22] ;
 wire \k[23] ;
 wire \k[24] ;
 wire \k[25] ;
 wire \k[26] ;
 wire \k[27] ;
 wire \k[28] ;
 wire \k[29] ;
 wire \k[2] ;
 wire \k[30] ;
 wire \k[31] ;
 wire \k[3] ;
 wire \k[4] ;
 wire \k[5] ;
 wire \k[6] ;
 wire \k[7] ;
 wire \k[8] ;
 wire \k[9] ;
 wire \second_row[0][0] ;
 wire \second_row[0][1] ;
 wire \second_row[0][2] ;
 wire \second_row[0][3] ;
 wire \second_row[0][4] ;
 wire \second_row[0][5] ;
 wire \second_row[0][6] ;
 wire \second_row[0][7] ;
 wire \second_row[10][0] ;
 wire \second_row[10][1] ;
 wire \second_row[10][2] ;
 wire \second_row[10][3] ;
 wire \second_row[10][4] ;
 wire \second_row[10][5] ;
 wire \second_row[10][6] ;
 wire \second_row[10][7] ;
 wire \second_row[11][0] ;
 wire \second_row[11][1] ;
 wire \second_row[11][2] ;
 wire \second_row[11][3] ;
 wire \second_row[11][4] ;
 wire \second_row[11][5] ;
 wire \second_row[11][6] ;
 wire \second_row[11][7] ;
 wire \second_row[12][0] ;
 wire \second_row[12][1] ;
 wire \second_row[12][2] ;
 wire \second_row[12][3] ;
 wire \second_row[12][4] ;
 wire \second_row[12][5] ;
 wire \second_row[12][6] ;
 wire \second_row[12][7] ;
 wire \second_row[13][0] ;
 wire \second_row[13][1] ;
 wire \second_row[13][2] ;
 wire \second_row[13][3] ;
 wire \second_row[13][4] ;
 wire \second_row[13][5] ;
 wire \second_row[13][6] ;
 wire \second_row[13][7] ;
 wire \second_row[14][0] ;
 wire \second_row[14][1] ;
 wire \second_row[14][2] ;
 wire \second_row[14][3] ;
 wire \second_row[14][4] ;
 wire \second_row[14][5] ;
 wire \second_row[14][6] ;
 wire \second_row[14][7] ;
 wire \second_row[15][0] ;
 wire \second_row[15][1] ;
 wire \second_row[15][2] ;
 wire \second_row[15][3] ;
 wire \second_row[15][4] ;
 wire \second_row[15][5] ;
 wire \second_row[15][6] ;
 wire \second_row[15][7] ;
 wire \second_row[16][0] ;
 wire \second_row[16][1] ;
 wire \second_row[16][2] ;
 wire \second_row[16][3] ;
 wire \second_row[16][4] ;
 wire \second_row[16][5] ;
 wire \second_row[16][6] ;
 wire \second_row[16][7] ;
 wire \second_row[17][0] ;
 wire \second_row[17][1] ;
 wire \second_row[17][2] ;
 wire \second_row[17][3] ;
 wire \second_row[17][4] ;
 wire \second_row[17][5] ;
 wire \second_row[17][6] ;
 wire \second_row[17][7] ;
 wire \second_row[1][0] ;
 wire \second_row[1][1] ;
 wire \second_row[1][2] ;
 wire \second_row[1][3] ;
 wire \second_row[1][4] ;
 wire \second_row[1][5] ;
 wire \second_row[1][6] ;
 wire \second_row[1][7] ;
 wire \second_row[2][0] ;
 wire \second_row[2][1] ;
 wire \second_row[2][2] ;
 wire \second_row[2][3] ;
 wire \second_row[2][4] ;
 wire \second_row[2][5] ;
 wire \second_row[2][6] ;
 wire \second_row[2][7] ;
 wire \second_row[3][0] ;
 wire \second_row[3][1] ;
 wire \second_row[3][2] ;
 wire \second_row[3][3] ;
 wire \second_row[3][4] ;
 wire \second_row[3][5] ;
 wire \second_row[3][6] ;
 wire \second_row[3][7] ;
 wire \second_row[4][0] ;
 wire \second_row[4][1] ;
 wire \second_row[4][2] ;
 wire \second_row[4][3] ;
 wire \second_row[4][4] ;
 wire \second_row[4][5] ;
 wire \second_row[4][6] ;
 wire \second_row[4][7] ;
 wire \second_row[5][0] ;
 wire \second_row[5][1] ;
 wire \second_row[5][2] ;
 wire \second_row[5][3] ;
 wire \second_row[5][4] ;
 wire \second_row[5][5] ;
 wire \second_row[5][6] ;
 wire \second_row[5][7] ;
 wire \second_row[6][0] ;
 wire \second_row[6][1] ;
 wire \second_row[6][2] ;
 wire \second_row[6][3] ;
 wire \second_row[6][4] ;
 wire \second_row[6][5] ;
 wire \second_row[6][6] ;
 wire \second_row[6][7] ;
 wire \second_row[7][0] ;
 wire \second_row[7][1] ;
 wire \second_row[7][2] ;
 wire \second_row[7][3] ;
 wire \second_row[7][4] ;
 wire \second_row[7][5] ;
 wire \second_row[7][6] ;
 wire \second_row[7][7] ;
 wire \second_row[8][0] ;
 wire \second_row[8][1] ;
 wire \second_row[8][2] ;
 wire \second_row[8][3] ;
 wire \second_row[8][4] ;
 wire \second_row[8][5] ;
 wire \second_row[8][6] ;
 wire \second_row[8][7] ;
 wire \second_row[9][0] ;
 wire \second_row[9][1] ;
 wire \second_row[9][2] ;
 wire \second_row[9][3] ;
 wire \second_row[9][4] ;
 wire \second_row[9][5] ;
 wire \second_row[9][6] ;
 wire \second_row[9][7] ;
 wire \third_row[0][0] ;
 wire \third_row[0][1] ;
 wire \third_row[0][2] ;
 wire \third_row[0][3] ;
 wire \third_row[0][4] ;
 wire \third_row[0][5] ;
 wire \third_row[0][6] ;
 wire \third_row[0][7] ;
 wire \third_row[10][0] ;
 wire \third_row[10][1] ;
 wire \third_row[10][2] ;
 wire \third_row[10][3] ;
 wire \third_row[10][4] ;
 wire \third_row[10][5] ;
 wire \third_row[10][6] ;
 wire \third_row[10][7] ;
 wire \third_row[11][0] ;
 wire \third_row[11][1] ;
 wire \third_row[11][2] ;
 wire \third_row[11][3] ;
 wire \third_row[11][4] ;
 wire \third_row[11][5] ;
 wire \third_row[11][6] ;
 wire \third_row[11][7] ;
 wire \third_row[12][0] ;
 wire \third_row[12][1] ;
 wire \third_row[12][2] ;
 wire \third_row[12][3] ;
 wire \third_row[12][4] ;
 wire \third_row[12][5] ;
 wire \third_row[12][6] ;
 wire \third_row[12][7] ;
 wire \third_row[13][0] ;
 wire \third_row[13][1] ;
 wire \third_row[13][2] ;
 wire \third_row[13][3] ;
 wire \third_row[13][4] ;
 wire \third_row[13][5] ;
 wire \third_row[13][6] ;
 wire \third_row[13][7] ;
 wire \third_row[14][0] ;
 wire \third_row[14][1] ;
 wire \third_row[14][2] ;
 wire \third_row[14][3] ;
 wire \third_row[14][4] ;
 wire \third_row[14][5] ;
 wire \third_row[14][6] ;
 wire \third_row[14][7] ;
 wire \third_row[15][0] ;
 wire \third_row[15][1] ;
 wire \third_row[15][2] ;
 wire \third_row[15][3] ;
 wire \third_row[15][4] ;
 wire \third_row[15][5] ;
 wire \third_row[15][6] ;
 wire \third_row[15][7] ;
 wire \third_row[16][0] ;
 wire \third_row[16][1] ;
 wire \third_row[16][2] ;
 wire \third_row[16][3] ;
 wire \third_row[16][4] ;
 wire \third_row[16][5] ;
 wire \third_row[16][6] ;
 wire \third_row[16][7] ;
 wire \third_row[17][0] ;
 wire \third_row[17][1] ;
 wire \third_row[17][2] ;
 wire \third_row[17][3] ;
 wire \third_row[17][4] ;
 wire \third_row[17][5] ;
 wire \third_row[17][6] ;
 wire \third_row[17][7] ;
 wire \third_row[1][0] ;
 wire \third_row[1][1] ;
 wire \third_row[1][2] ;
 wire \third_row[1][3] ;
 wire \third_row[1][4] ;
 wire \third_row[1][5] ;
 wire \third_row[1][6] ;
 wire \third_row[1][7] ;
 wire \third_row[2][0] ;
 wire \third_row[2][1] ;
 wire \third_row[2][2] ;
 wire \third_row[2][3] ;
 wire \third_row[2][4] ;
 wire \third_row[2][5] ;
 wire \third_row[2][6] ;
 wire \third_row[2][7] ;
 wire \third_row[3][0] ;
 wire \third_row[3][1] ;
 wire \third_row[3][2] ;
 wire \third_row[3][3] ;
 wire \third_row[3][4] ;
 wire \third_row[3][5] ;
 wire \third_row[3][6] ;
 wire \third_row[3][7] ;
 wire \third_row[4][0] ;
 wire \third_row[4][1] ;
 wire \third_row[4][2] ;
 wire \third_row[4][3] ;
 wire \third_row[4][4] ;
 wire \third_row[4][5] ;
 wire \third_row[4][6] ;
 wire \third_row[4][7] ;
 wire \third_row[5][0] ;
 wire \third_row[5][1] ;
 wire \third_row[5][2] ;
 wire \third_row[5][3] ;
 wire \third_row[5][4] ;
 wire \third_row[5][5] ;
 wire \third_row[5][6] ;
 wire \third_row[5][7] ;
 wire \third_row[6][0] ;
 wire \third_row[6][1] ;
 wire \third_row[6][2] ;
 wire \third_row[6][3] ;
 wire \third_row[6][4] ;
 wire \third_row[6][5] ;
 wire \third_row[6][6] ;
 wire \third_row[6][7] ;
 wire \third_row[7][0] ;
 wire \third_row[7][1] ;
 wire \third_row[7][2] ;
 wire \third_row[7][3] ;
 wire \third_row[7][4] ;
 wire \third_row[7][5] ;
 wire \third_row[7][6] ;
 wire \third_row[7][7] ;
 wire \third_row[8][0] ;
 wire \third_row[8][1] ;
 wire \third_row[8][2] ;
 wire \third_row[8][3] ;
 wire \third_row[8][4] ;
 wire \third_row[8][5] ;
 wire \third_row[8][6] ;
 wire \third_row[8][7] ;
 wire \third_row[9][0] ;
 wire \third_row[9][1] ;
 wire \third_row[9][2] ;
 wire \third_row[9][3] ;
 wire \third_row[9][4] ;
 wire \third_row[9][5] ;
 wire \third_row[9][6] ;
 wire \third_row[9][7] ;
 wire \valid_counter[0] ;
 wire \valid_counter[10] ;
 wire \valid_counter[11] ;
 wire \valid_counter[12] ;
 wire \valid_counter[13] ;
 wire \valid_counter[14] ;
 wire \valid_counter[15] ;
 wire \valid_counter[16] ;
 wire \valid_counter[17] ;
 wire \valid_counter[18] ;
 wire \valid_counter[19] ;
 wire \valid_counter[1] ;
 wire \valid_counter[20] ;
 wire \valid_counter[21] ;
 wire \valid_counter[22] ;
 wire \valid_counter[23] ;
 wire \valid_counter[24] ;
 wire \valid_counter[25] ;
 wire \valid_counter[26] ;
 wire \valid_counter[27] ;
 wire \valid_counter[28] ;
 wire \valid_counter[29] ;
 wire \valid_counter[2] ;
 wire \valid_counter[30] ;
 wire \valid_counter[31] ;
 wire \valid_counter[3] ;
 wire \valid_counter[4] ;
 wire \valid_counter[5] ;
 wire \valid_counter[6] ;
 wire \valid_counter[7] ;
 wire \valid_counter[8] ;
 wire \valid_counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_leaf_0_CLK;
 wire clknet_leaf_1_CLK;
 wire clknet_leaf_2_CLK;
 wire clknet_leaf_3_CLK;
 wire clknet_leaf_4_CLK;
 wire clknet_leaf_5_CLK;
 wire clknet_leaf_6_CLK;
 wire clknet_leaf_7_CLK;
 wire clknet_leaf_8_CLK;
 wire clknet_leaf_9_CLK;
 wire clknet_leaf_10_CLK;
 wire clknet_leaf_11_CLK;
 wire clknet_leaf_12_CLK;
 wire clknet_leaf_13_CLK;
 wire clknet_leaf_14_CLK;
 wire clknet_leaf_15_CLK;
 wire clknet_leaf_16_CLK;
 wire clknet_leaf_17_CLK;
 wire clknet_leaf_18_CLK;
 wire clknet_leaf_19_CLK;
 wire clknet_leaf_20_CLK;
 wire clknet_leaf_21_CLK;
 wire clknet_leaf_22_CLK;
 wire clknet_leaf_23_CLK;
 wire clknet_leaf_24_CLK;
 wire clknet_leaf_25_CLK;
 wire clknet_leaf_26_CLK;
 wire clknet_leaf_28_CLK;
 wire clknet_leaf_29_CLK;
 wire clknet_leaf_30_CLK;
 wire clknet_leaf_31_CLK;
 wire clknet_leaf_32_CLK;
 wire clknet_leaf_33_CLK;
 wire clknet_leaf_34_CLK;
 wire clknet_leaf_35_CLK;
 wire clknet_leaf_36_CLK;
 wire clknet_leaf_37_CLK;
 wire clknet_leaf_38_CLK;
 wire clknet_leaf_39_CLK;
 wire clknet_leaf_40_CLK;
 wire clknet_leaf_41_CLK;
 wire clknet_leaf_42_CLK;
 wire clknet_leaf_43_CLK;
 wire clknet_leaf_44_CLK;
 wire clknet_leaf_45_CLK;
 wire clknet_leaf_46_CLK;
 wire clknet_leaf_47_CLK;
 wire clknet_leaf_48_CLK;
 wire clknet_leaf_49_CLK;
 wire clknet_leaf_50_CLK;
 wire clknet_leaf_51_CLK;
 wire clknet_leaf_52_CLK;
 wire clknet_leaf_53_CLK;
 wire clknet_leaf_54_CLK;
 wire clknet_leaf_55_CLK;
 wire clknet_leaf_56_CLK;
 wire clknet_leaf_57_CLK;
 wire clknet_leaf_58_CLK;
 wire clknet_leaf_59_CLK;
 wire clknet_leaf_60_CLK;
 wire clknet_leaf_61_CLK;
 wire clknet_leaf_62_CLK;
 wire clknet_leaf_63_CLK;
 wire clknet_leaf_64_CLK;
 wire clknet_0_CLK;
 wire clknet_3_0__leaf_CLK;
 wire clknet_3_1__leaf_CLK;
 wire clknet_3_2__leaf_CLK;
 wire clknet_3_3__leaf_CLK;
 wire clknet_3_4__leaf_CLK;
 wire clknet_3_5__leaf_CLK;
 wire clknet_3_6__leaf_CLK;
 wire clknet_3_7__leaf_CLK;

 sky130_fd_sc_hd__inv_2 _2607_ (.A(net10),
    .Y(_1067_));
 sky130_fd_sc_hd__or4_1 _2608_ (.A(\col_input[11] ),
    .B(\col_input[10] ),
    .C(\col_input[9] ),
    .D(\col_input[8] ),
    .X(_1068_));
 sky130_fd_sc_hd__or3_1 _2609_ (.A(\col_input[15] ),
    .B(\col_input[14] ),
    .C(\col_input[13] ),
    .X(_1069_));
 sky130_fd_sc_hd__or4_1 _2610_ (.A(\col_input[12] ),
    .B(\col_input[7] ),
    .C(\col_input[6] ),
    .D(\col_input[5] ),
    .X(_1070_));
 sky130_fd_sc_hd__or3_1 _2611_ (.A(_1068_),
    .B(_1069_),
    .C(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__or4_1 _2612_ (.A(\col_input[27] ),
    .B(\col_input[26] ),
    .C(\col_input[25] ),
    .D(\col_input[24] ),
    .X(_1072_));
 sky130_fd_sc_hd__or4_1 _2613_ (.A(\col_input[31] ),
    .B(\col_input[30] ),
    .C(\col_input[29] ),
    .D(\col_input[28] ),
    .X(_1073_));
 sky130_fd_sc_hd__or4_1 _2614_ (.A(\col_input[19] ),
    .B(\col_input[18] ),
    .C(\col_input[17] ),
    .D(\col_input[16] ),
    .X(_1074_));
 sky130_fd_sc_hd__or4_1 _2615_ (.A(\col_input[23] ),
    .B(\col_input[22] ),
    .C(\col_input[21] ),
    .D(\col_input[20] ),
    .X(_1075_));
 sky130_fd_sc_hd__or4_2 _2616_ (.A(_1072_),
    .B(_1073_),
    .C(_1074_),
    .D(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__buf_2 _2617_ (.A(\col_input[3] ),
    .X(_1077_));
 sky130_fd_sc_hd__or4b_1 _2618_ (.A(_1077_),
    .B(\col_input[2] ),
    .C(\col_input[1] ),
    .D_N(\col_input[0] ),
    .X(_1078_));
 sky130_fd_sc_hd__or4_2 _2619_ (.A(\col_input[4] ),
    .B(_1071_),
    .C(_1076_),
    .D(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__or2_1 _2620_ (.A(_1067_),
    .B(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_4 _2621_ (.A(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__clkbuf_8 _2622_ (.A(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__buf_4 _2623_ (.A(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(\second_row[17][7] ),
    .A1(\third_row[17][7] ),
    .S(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2625_ (.A(_1084_),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(\second_row[17][6] ),
    .A1(\third_row[17][6] ),
    .S(_1083_),
    .X(_1085_));
 sky130_fd_sc_hd__clkbuf_1 _2627_ (.A(_1085_),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(\second_row[17][5] ),
    .A1(\third_row[17][5] ),
    .S(_1083_),
    .X(_1086_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_1086_),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(\second_row[17][4] ),
    .A1(\third_row[17][4] ),
    .S(_1083_),
    .X(_1087_));
 sky130_fd_sc_hd__clkbuf_1 _2631_ (.A(_1087_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(\second_row[17][3] ),
    .A1(\third_row[17][3] ),
    .S(_1083_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_1 _2633_ (.A(_1088_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\second_row[17][2] ),
    .A1(\third_row[17][2] ),
    .S(_1083_),
    .X(_1089_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1089_),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(\second_row[17][1] ),
    .A1(\third_row[17][1] ),
    .S(_1083_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_1090_),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(\second_row[17][0] ),
    .A1(\third_row[17][0] ),
    .S(_1083_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_1091_),
    .X(_1059_));
 sky130_fd_sc_hd__buf_2 _2640_ (.A(net8),
    .X(_1092_));
 sky130_fd_sc_hd__nor2_2 _2641_ (.A(\col_input[3] ),
    .B(\col_input[2] ),
    .Y(_1093_));
 sky130_fd_sc_hd__inv_2 _2642_ (.A(\col_input[4] ),
    .Y(_1094_));
 sky130_fd_sc_hd__nor2_1 _2643_ (.A(\col_input[1] ),
    .B(\col_input[0] ),
    .Y(_1095_));
 sky130_fd_sc_hd__a21oi_1 _2644_ (.A1(_1093_),
    .A2(_1095_),
    .B1(_1094_),
    .Y(_1096_));
 sky130_fd_sc_hd__inv_2 _2645_ (.A(\col_input[31] ),
    .Y(_1097_));
 sky130_fd_sc_hd__o31a_1 _2646_ (.A1(_1071_),
    .A2(_1076_),
    .A3(_1096_),
    .B1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__nor2_2 _2647_ (.A(_1067_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__and3_4 _2648_ (.A(_1094_),
    .B(_1095_),
    .C(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__nand2_4 _2649_ (.A(_1093_),
    .B(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(_1092_),
    .A1(\first_row[0][7] ),
    .S(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_1102_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_2 _2652_ (.A(net7),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(_1103_),
    .A1(\first_row[0][6] ),
    .S(_1101_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2654_ (.A(_1104_),
    .X(_1057_));
 sky130_fd_sc_hd__buf_2 _2655_ (.A(net6),
    .X(_1105_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(_1105_),
    .A1(\first_row[0][5] ),
    .S(_1101_),
    .X(_1106_));
 sky130_fd_sc_hd__clkbuf_1 _2657_ (.A(_1106_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_2 _2658_ (.A(net5),
    .X(_1107_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(_1107_),
    .A1(\first_row[0][4] ),
    .S(_1101_),
    .X(_1108_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1108_),
    .X(_1055_));
 sky130_fd_sc_hd__clkbuf_2 _2661_ (.A(net4),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(_1109_),
    .A1(\first_row[0][3] ),
    .S(_1101_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(_1110_),
    .X(_1054_));
 sky130_fd_sc_hd__clkbuf_2 _2664_ (.A(net3),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(_1111_),
    .A1(\first_row[0][2] ),
    .S(_1101_),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_1112_),
    .X(_1053_));
 sky130_fd_sc_hd__clkbuf_2 _2667_ (.A(net2),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(_1113_),
    .A1(\first_row[0][1] ),
    .S(_1101_),
    .X(_1114_));
 sky130_fd_sc_hd__clkbuf_1 _2669_ (.A(_1114_),
    .X(_1052_));
 sky130_fd_sc_hd__buf_2 _2670_ (.A(net1),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _2671_ (.A0(_1115_),
    .A1(\first_row[0][0] ),
    .S(_1101_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_1116_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2673_ (.A0(\second_row[16][7] ),
    .A1(\third_row[16][7] ),
    .S(_1083_),
    .X(_1117_));
 sky130_fd_sc_hd__clkbuf_1 _2674_ (.A(_1117_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(\second_row[16][6] ),
    .A1(\third_row[16][6] ),
    .S(_1083_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _2676_ (.A(_1118_),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_8 _2677_ (.A(_1082_),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(\second_row[16][5] ),
    .A1(\third_row[16][5] ),
    .S(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _2679_ (.A(_1120_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(\second_row[16][4] ),
    .A1(\third_row[16][4] ),
    .S(_1119_),
    .X(_1121_));
 sky130_fd_sc_hd__clkbuf_1 _2681_ (.A(_1121_),
    .X(_1047_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(\second_row[16][3] ),
    .A1(\third_row[16][3] ),
    .S(_1119_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2683_ (.A(_1122_),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(\second_row[16][2] ),
    .A1(\third_row[16][2] ),
    .S(_1119_),
    .X(_1123_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1123_),
    .X(_1045_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(\second_row[16][1] ),
    .A1(\third_row[16][1] ),
    .S(_1119_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_1 _2687_ (.A(_1124_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(\second_row[16][0] ),
    .A1(\third_row[16][0] ),
    .S(_1119_),
    .X(_1125_));
 sky130_fd_sc_hd__clkbuf_1 _2689_ (.A(_1125_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(\second_row[15][7] ),
    .A1(\third_row[15][7] ),
    .S(_1119_),
    .X(_1126_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1126_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(\second_row[15][6] ),
    .A1(\third_row[15][6] ),
    .S(_1119_),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1127_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\second_row[15][5] ),
    .A1(\third_row[15][5] ),
    .S(_1119_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1128_),
    .X(_1040_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(\second_row[15][4] ),
    .A1(\third_row[15][4] ),
    .S(_1119_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1129_),
    .X(_1039_));
 sky130_fd_sc_hd__buf_2 _2698_ (.A(_1081_),
    .X(_1130_));
 sky130_fd_sc_hd__buf_4 _2699_ (.A(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(\second_row[15][3] ),
    .A1(\third_row[15][3] ),
    .S(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2701_ (.A(_1132_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(\second_row[15][2] ),
    .A1(\third_row[15][2] ),
    .S(_1131_),
    .X(_1133_));
 sky130_fd_sc_hd__clkbuf_1 _2703_ (.A(_1133_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(\second_row[15][1] ),
    .A1(\third_row[15][1] ),
    .S(_1131_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2705_ (.A(_1134_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _2706_ (.A0(\second_row[15][0] ),
    .A1(\third_row[15][0] ),
    .S(_1131_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2707_ (.A(_1135_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2708_ (.A0(\second_row[14][7] ),
    .A1(\third_row[14][7] ),
    .S(_1131_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _2709_ (.A(_1136_),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\second_row[14][6] ),
    .A1(\third_row[14][6] ),
    .S(_1131_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _2711_ (.A(_1137_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _2712_ (.A0(\second_row[14][5] ),
    .A1(\third_row[14][5] ),
    .S(_1131_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_1 _2713_ (.A(_1138_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(\second_row[14][4] ),
    .A1(\third_row[14][4] ),
    .S(_1131_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _2715_ (.A(_1139_),
    .X(_1031_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\second_row[14][3] ),
    .A1(\third_row[14][3] ),
    .S(_1131_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _2717_ (.A(_1140_),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(\second_row[14][2] ),
    .A1(\third_row[14][2] ),
    .S(_1131_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2719_ (.A(_1141_),
    .X(_1029_));
 sky130_fd_sc_hd__buf_4 _2720_ (.A(_1130_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(\second_row[14][1] ),
    .A1(\third_row[14][1] ),
    .S(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _2722_ (.A(_1143_),
    .X(_1028_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(\second_row[14][0] ),
    .A1(\third_row[14][0] ),
    .S(_1142_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2724_ (.A(_1144_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _2725_ (.A0(\second_row[13][7] ),
    .A1(\third_row[13][7] ),
    .S(_1142_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _2726_ (.A(_1145_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(\second_row[13][6] ),
    .A1(\third_row[13][6] ),
    .S(_1142_),
    .X(_1146_));
 sky130_fd_sc_hd__clkbuf_1 _2728_ (.A(_1146_),
    .X(_1025_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(\second_row[13][5] ),
    .A1(\third_row[13][5] ),
    .S(_1142_),
    .X(_1147_));
 sky130_fd_sc_hd__clkbuf_1 _2730_ (.A(_1147_),
    .X(_1024_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(\second_row[13][4] ),
    .A1(\third_row[13][4] ),
    .S(_1142_),
    .X(_1148_));
 sky130_fd_sc_hd__clkbuf_1 _2732_ (.A(_1148_),
    .X(_1023_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(\second_row[13][3] ),
    .A1(\third_row[13][3] ),
    .S(_1142_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_1 _2734_ (.A(_1149_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(\second_row[13][2] ),
    .A1(\third_row[13][2] ),
    .S(_1142_),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2736_ (.A(_1150_),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(\second_row[13][1] ),
    .A1(\third_row[13][1] ),
    .S(_1142_),
    .X(_1151_));
 sky130_fd_sc_hd__clkbuf_1 _2738_ (.A(_1151_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(\second_row[13][0] ),
    .A1(\third_row[13][0] ),
    .S(_1142_),
    .X(_1152_));
 sky130_fd_sc_hd__clkbuf_1 _2740_ (.A(_1152_),
    .X(_1019_));
 sky130_fd_sc_hd__buf_4 _2741_ (.A(_1130_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(\second_row[12][7] ),
    .A1(\third_row[12][7] ),
    .S(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__clkbuf_1 _2743_ (.A(_1154_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(\second_row[12][6] ),
    .A1(\third_row[12][6] ),
    .S(_1153_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1155_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(\second_row[12][5] ),
    .A1(\third_row[12][5] ),
    .S(_1153_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2747_ (.A(_1156_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\second_row[12][4] ),
    .A1(\third_row[12][4] ),
    .S(_1153_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2749_ (.A(_1157_),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(\second_row[12][3] ),
    .A1(\third_row[12][3] ),
    .S(_1153_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_1 _2751_ (.A(_1158_),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(\second_row[12][2] ),
    .A1(\third_row[12][2] ),
    .S(_1153_),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _2753_ (.A(_1159_),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(\second_row[12][1] ),
    .A1(\third_row[12][1] ),
    .S(_1153_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_1 _2755_ (.A(_1160_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _2756_ (.A0(\second_row[12][0] ),
    .A1(\third_row[12][0] ),
    .S(_1153_),
    .X(_1161_));
 sky130_fd_sc_hd__clkbuf_1 _2757_ (.A(_1161_),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _2758_ (.A0(\second_row[11][7] ),
    .A1(\third_row[11][7] ),
    .S(_1153_),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _2759_ (.A(_1162_),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(\second_row[11][6] ),
    .A1(\third_row[11][6] ),
    .S(_1153_),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_1 _2761_ (.A(_1163_),
    .X(_1009_));
 sky130_fd_sc_hd__buf_4 _2762_ (.A(_1130_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(\second_row[11][5] ),
    .A1(\third_row[11][5] ),
    .S(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_1165_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(\second_row[11][4] ),
    .A1(\third_row[11][4] ),
    .S(_1164_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(_1166_),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(\second_row[11][3] ),
    .A1(\third_row[11][3] ),
    .S(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(_1167_),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(\second_row[11][2] ),
    .A1(\third_row[11][2] ),
    .S(_1164_),
    .X(_1168_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_1168_),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(\second_row[11][1] ),
    .A1(\third_row[11][1] ),
    .S(_1164_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _2772_ (.A(_1169_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(\second_row[11][0] ),
    .A1(\third_row[11][0] ),
    .S(_1164_),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _2774_ (.A(_1170_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\second_row[10][7] ),
    .A1(\third_row[10][7] ),
    .S(_1164_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _2776_ (.A(_1171_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\second_row[10][6] ),
    .A1(\third_row[10][6] ),
    .S(_1164_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _2778_ (.A(_1172_),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\second_row[10][5] ),
    .A1(\third_row[10][5] ),
    .S(_1164_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2780_ (.A(_1173_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\second_row[10][4] ),
    .A1(\third_row[10][4] ),
    .S(_1164_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2782_ (.A(_1174_),
    .X(_0999_));
 sky130_fd_sc_hd__buf_4 _2783_ (.A(_1130_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(\second_row[10][3] ),
    .A1(\third_row[10][3] ),
    .S(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__clkbuf_1 _2785_ (.A(_1176_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(\second_row[10][2] ),
    .A1(\third_row[10][2] ),
    .S(_1175_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _2787_ (.A(_1177_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(\second_row[10][1] ),
    .A1(\third_row[10][1] ),
    .S(_1175_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2789_ (.A(_1178_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\second_row[10][0] ),
    .A1(\third_row[10][0] ),
    .S(_1175_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2791_ (.A(_1179_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\second_row[9][7] ),
    .A1(\third_row[9][7] ),
    .S(_1175_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2793_ (.A(_1180_),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\second_row[9][6] ),
    .A1(\third_row[9][6] ),
    .S(_1175_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _2795_ (.A(_1181_),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\second_row[9][5] ),
    .A1(\third_row[9][5] ),
    .S(_1175_),
    .X(_1182_));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(_1182_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\second_row[9][4] ),
    .A1(\third_row[9][4] ),
    .S(_1175_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _2799_ (.A(_1183_),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\second_row[9][3] ),
    .A1(\third_row[9][3] ),
    .S(_1175_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(_1184_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\second_row[9][2] ),
    .A1(\third_row[9][2] ),
    .S(_1175_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1185_),
    .X(_0989_));
 sky130_fd_sc_hd__buf_4 _2804_ (.A(_1130_),
    .X(_1186_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\second_row[9][1] ),
    .A1(\third_row[9][1] ),
    .S(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _2806_ (.A(_1187_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(\second_row[9][0] ),
    .A1(\third_row[9][0] ),
    .S(_1186_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2808_ (.A(_1188_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\second_row[8][7] ),
    .A1(\third_row[8][7] ),
    .S(_1186_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2810_ (.A(_1189_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(\second_row[8][6] ),
    .A1(\third_row[8][6] ),
    .S(_1186_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2812_ (.A(_1190_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(\second_row[8][5] ),
    .A1(\third_row[8][5] ),
    .S(_1186_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2814_ (.A(_1191_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(\second_row[8][4] ),
    .A1(\third_row[8][4] ),
    .S(_1186_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _2816_ (.A(_1192_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(\second_row[8][3] ),
    .A1(\third_row[8][3] ),
    .S(_1186_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2818_ (.A(_1193_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(\second_row[8][2] ),
    .A1(\third_row[8][2] ),
    .S(_1186_),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_1 _2820_ (.A(_1194_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(\second_row[8][1] ),
    .A1(\third_row[8][1] ),
    .S(_1186_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2822_ (.A(_1195_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(\second_row[8][0] ),
    .A1(\third_row[8][0] ),
    .S(_1186_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2824_ (.A(_1196_),
    .X(_0979_));
 sky130_fd_sc_hd__buf_4 _2825_ (.A(_1130_),
    .X(_1197_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(\second_row[7][7] ),
    .A1(\third_row[7][7] ),
    .S(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2827_ (.A(_1198_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(\second_row[7][6] ),
    .A1(\third_row[7][6] ),
    .S(_1197_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2829_ (.A(_1199_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(\second_row[7][5] ),
    .A1(\third_row[7][5] ),
    .S(_1197_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _2831_ (.A(_1200_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(\second_row[7][4] ),
    .A1(\third_row[7][4] ),
    .S(_1197_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2833_ (.A(_1201_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _2834_ (.A0(\second_row[7][3] ),
    .A1(\third_row[7][3] ),
    .S(_1197_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2835_ (.A(_1202_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(\second_row[7][2] ),
    .A1(\third_row[7][2] ),
    .S(_1197_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2837_ (.A(_1203_),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(\second_row[7][1] ),
    .A1(\third_row[7][1] ),
    .S(_1197_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2839_ (.A(_1204_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(\second_row[7][0] ),
    .A1(\third_row[7][0] ),
    .S(_1197_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2841_ (.A(_1205_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(\second_row[6][7] ),
    .A1(\third_row[6][7] ),
    .S(_1197_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2843_ (.A(_1206_),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(\second_row[6][6] ),
    .A1(\third_row[6][6] ),
    .S(_1197_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_1207_),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_4 _2846_ (.A(_1130_),
    .X(_1208_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(\second_row[6][5] ),
    .A1(\third_row[6][5] ),
    .S(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2848_ (.A(_1209_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(\second_row[6][4] ),
    .A1(\third_row[6][4] ),
    .S(_1208_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1210_),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\second_row[6][3] ),
    .A1(\third_row[6][3] ),
    .S(_1208_),
    .X(_1211_));
 sky130_fd_sc_hd__clkbuf_1 _2852_ (.A(_1211_),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\second_row[6][2] ),
    .A1(\third_row[6][2] ),
    .S(_1208_),
    .X(_1212_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1212_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\second_row[6][1] ),
    .A1(\third_row[6][1] ),
    .S(_1208_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2856_ (.A(_1213_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\second_row[6][0] ),
    .A1(\third_row[6][0] ),
    .S(_1208_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _2858_ (.A(_1214_),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\second_row[5][7] ),
    .A1(\third_row[5][7] ),
    .S(_1208_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(_1215_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(\second_row[5][6] ),
    .A1(\third_row[5][6] ),
    .S(_1208_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _2862_ (.A(_1216_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(\second_row[5][5] ),
    .A1(\third_row[5][5] ),
    .S(_1208_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _2864_ (.A(_1217_),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\second_row[5][4] ),
    .A1(\third_row[5][4] ),
    .S(_1208_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1218_),
    .X(_0959_));
 sky130_fd_sc_hd__buf_4 _2867_ (.A(_1130_),
    .X(_1219_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\second_row[5][3] ),
    .A1(\third_row[5][3] ),
    .S(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_1220_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\second_row[5][2] ),
    .A1(\third_row[5][2] ),
    .S(_1219_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2871_ (.A(_1221_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\second_row[5][1] ),
    .A1(\third_row[5][1] ),
    .S(_1219_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2873_ (.A(_1222_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\second_row[5][0] ),
    .A1(\third_row[5][0] ),
    .S(_1219_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1223_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\second_row[4][7] ),
    .A1(\third_row[4][7] ),
    .S(_1219_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1224_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(\second_row[4][6] ),
    .A1(\third_row[4][6] ),
    .S(_1219_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_1225_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(\second_row[4][5] ),
    .A1(\third_row[4][5] ),
    .S(_1219_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2881_ (.A(_1226_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(\second_row[4][4] ),
    .A1(\third_row[4][4] ),
    .S(_1219_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2883_ (.A(_1227_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(\second_row[4][3] ),
    .A1(\third_row[4][3] ),
    .S(_1219_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(_1228_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(\second_row[4][2] ),
    .A1(\third_row[4][2] ),
    .S(_1219_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2887_ (.A(_1229_),
    .X(_0949_));
 sky130_fd_sc_hd__buf_4 _2888_ (.A(_1130_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(\second_row[4][1] ),
    .A1(\third_row[4][1] ),
    .S(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2890_ (.A(_1231_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(\second_row[4][0] ),
    .A1(\third_row[4][0] ),
    .S(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1232_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(\second_row[3][7] ),
    .A1(\third_row[3][7] ),
    .S(_1230_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2894_ (.A(_1233_),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(\second_row[3][6] ),
    .A1(\third_row[3][6] ),
    .S(_1230_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2896_ (.A(_1234_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(\second_row[3][5] ),
    .A1(\third_row[3][5] ),
    .S(_1230_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_1235_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(\second_row[3][4] ),
    .A1(\third_row[3][4] ),
    .S(_1230_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2900_ (.A(_1236_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(\second_row[3][3] ),
    .A1(\third_row[3][3] ),
    .S(_1230_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2902_ (.A(_1237_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(\second_row[3][2] ),
    .A1(\third_row[3][2] ),
    .S(_1230_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2904_ (.A(_1238_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(\second_row[3][1] ),
    .A1(\third_row[3][1] ),
    .S(_1230_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _2906_ (.A(_1239_),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(\second_row[3][0] ),
    .A1(\third_row[3][0] ),
    .S(_1230_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1240_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_4 _2909_ (.A(_1081_),
    .X(_1241_));
 sky130_fd_sc_hd__buf_4 _2910_ (.A(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(\second_row[2][7] ),
    .A1(\third_row[2][7] ),
    .S(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1243_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(\second_row[2][6] ),
    .A1(\third_row[2][6] ),
    .S(_1242_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1244_),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(\second_row[2][5] ),
    .A1(\third_row[2][5] ),
    .S(_1242_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2916_ (.A(_1245_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(\second_row[2][4] ),
    .A1(\third_row[2][4] ),
    .S(_1242_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2918_ (.A(_1246_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(\second_row[2][3] ),
    .A1(\third_row[2][3] ),
    .S(_1242_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _2920_ (.A(_1247_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(\second_row[2][2] ),
    .A1(\third_row[2][2] ),
    .S(_1242_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _2922_ (.A(_1248_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(\second_row[2][1] ),
    .A1(\third_row[2][1] ),
    .S(_1242_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2924_ (.A(_1249_),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(\second_row[2][0] ),
    .A1(\third_row[2][0] ),
    .S(_1242_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2926_ (.A(_1250_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(\second_row[1][7] ),
    .A1(\third_row[1][7] ),
    .S(_1242_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2928_ (.A(_1251_),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(\second_row[1][6] ),
    .A1(\third_row[1][6] ),
    .S(_1242_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1252_),
    .X(_0929_));
 sky130_fd_sc_hd__clkbuf_8 _2931_ (.A(_1241_),
    .X(_1253_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(\second_row[1][5] ),
    .A1(\third_row[1][5] ),
    .S(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2933_ (.A(_1254_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(\second_row[1][4] ),
    .A1(\third_row[1][4] ),
    .S(_1253_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2935_ (.A(_1255_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _2936_ (.A0(\second_row[1][3] ),
    .A1(\third_row[1][3] ),
    .S(_1253_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2937_ (.A(_1256_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(\second_row[1][2] ),
    .A1(\third_row[1][2] ),
    .S(_1253_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1257_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(\second_row[1][1] ),
    .A1(\third_row[1][1] ),
    .S(_1253_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1258_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(\second_row[1][0] ),
    .A1(\third_row[1][0] ),
    .S(_1253_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2943_ (.A(_1259_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _2944_ (.A0(\second_row[0][7] ),
    .A1(\third_row[0][7] ),
    .S(_1253_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_1260_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(\second_row[0][6] ),
    .A1(\third_row[0][6] ),
    .S(_1253_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2947_ (.A(_1261_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(\second_row[0][5] ),
    .A1(\third_row[0][5] ),
    .S(_1253_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _2949_ (.A(_1262_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(\second_row[0][4] ),
    .A1(\third_row[0][4] ),
    .S(_1253_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2951_ (.A(_1263_),
    .X(_0919_));
 sky130_fd_sc_hd__buf_4 _2952_ (.A(_1241_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(\second_row[0][3] ),
    .A1(\third_row[0][3] ),
    .S(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1265_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(\second_row[0][2] ),
    .A1(\third_row[0][2] ),
    .S(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1266_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(\second_row[0][1] ),
    .A1(\third_row[0][1] ),
    .S(_1264_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1267_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(\second_row[0][0] ),
    .A1(\third_row[0][0] ),
    .S(_1264_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2960_ (.A(_1268_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(\first_row[17][7] ),
    .A1(\second_row[17][7] ),
    .S(_1264_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_1269_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(\first_row[17][6] ),
    .A1(\second_row[17][6] ),
    .S(_1264_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _2964_ (.A(_1270_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(\first_row[17][5] ),
    .A1(\second_row[17][5] ),
    .S(_1264_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_1271_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(\first_row[17][4] ),
    .A1(\second_row[17][4] ),
    .S(_1264_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1272_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(\first_row[17][3] ),
    .A1(\second_row[17][3] ),
    .S(_1264_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1273_),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(\first_row[17][2] ),
    .A1(\second_row[17][2] ),
    .S(_1264_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1274_),
    .X(_0909_));
 sky130_fd_sc_hd__buf_4 _2973_ (.A(_1241_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(\first_row[17][1] ),
    .A1(\second_row[17][1] ),
    .S(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2975_ (.A(_1276_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(\first_row[17][0] ),
    .A1(\second_row[17][0] ),
    .S(_1275_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1277_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(\first_row[16][7] ),
    .A1(\second_row[16][7] ),
    .S(_1275_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1278_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\first_row[16][6] ),
    .A1(\second_row[16][6] ),
    .S(_1275_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1279_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\first_row[16][5] ),
    .A1(\second_row[16][5] ),
    .S(_1275_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1280_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(\first_row[16][4] ),
    .A1(\second_row[16][4] ),
    .S(_1275_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2985_ (.A(_1281_),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(\first_row[16][3] ),
    .A1(\second_row[16][3] ),
    .S(_1275_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2987_ (.A(_1282_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(\first_row[16][2] ),
    .A1(\second_row[16][2] ),
    .S(_1275_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _2989_ (.A(_1283_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(\first_row[16][1] ),
    .A1(\second_row[16][1] ),
    .S(_1275_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2991_ (.A(_1284_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(\first_row[16][0] ),
    .A1(\second_row[16][0] ),
    .S(_1275_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _2993_ (.A(_1285_),
    .X(_0899_));
 sky130_fd_sc_hd__buf_4 _2994_ (.A(_1241_),
    .X(_1286_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(\first_row[15][7] ),
    .A1(\second_row[15][7] ),
    .S(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2996_ (.A(_1287_),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(\first_row[15][6] ),
    .A1(\second_row[15][6] ),
    .S(_1286_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_1288_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(\first_row[15][5] ),
    .A1(\second_row[15][5] ),
    .S(_1286_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _3000_ (.A(_1289_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(\first_row[15][4] ),
    .A1(\second_row[15][4] ),
    .S(_1286_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_1290_),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(\first_row[15][3] ),
    .A1(\second_row[15][3] ),
    .S(_1286_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _3004_ (.A(_1291_),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(\first_row[15][2] ),
    .A1(\second_row[15][2] ),
    .S(_1286_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1292_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(\first_row[15][1] ),
    .A1(\second_row[15][1] ),
    .S(_1286_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _3008_ (.A(_1293_),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(\first_row[15][0] ),
    .A1(\second_row[15][0] ),
    .S(_1286_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _3010_ (.A(_1294_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(\first_row[14][7] ),
    .A1(\second_row[14][7] ),
    .S(_1286_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _3012_ (.A(_1295_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(\first_row[14][6] ),
    .A1(\second_row[14][6] ),
    .S(_1286_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _3014_ (.A(_1296_),
    .X(_0889_));
 sky130_fd_sc_hd__buf_4 _3015_ (.A(_1241_),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(\first_row[14][5] ),
    .A1(\second_row[14][5] ),
    .S(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_1298_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\first_row[14][4] ),
    .A1(\second_row[14][4] ),
    .S(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1299_),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(\first_row[14][3] ),
    .A1(\second_row[14][3] ),
    .S(_1297_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1300_),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(\first_row[14][2] ),
    .A1(\second_row[14][2] ),
    .S(_1297_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1301_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(\first_row[14][1] ),
    .A1(\second_row[14][1] ),
    .S(_1297_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1302_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(\first_row[14][0] ),
    .A1(\second_row[14][0] ),
    .S(_1297_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_1303_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(\first_row[13][7] ),
    .A1(\second_row[13][7] ),
    .S(_1297_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _3029_ (.A(_1304_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(\first_row[13][6] ),
    .A1(\second_row[13][6] ),
    .S(_1297_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_1305_),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(\first_row[13][5] ),
    .A1(\second_row[13][5] ),
    .S(_1297_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1306_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(\first_row[13][4] ),
    .A1(\second_row[13][4] ),
    .S(_1297_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1307_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_8 _3036_ (.A(_1241_),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(\first_row[13][3] ),
    .A1(\second_row[13][3] ),
    .S(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _3038_ (.A(_1309_),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(\first_row[13][2] ),
    .A1(\second_row[13][2] ),
    .S(_1308_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _3040_ (.A(_1310_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(\first_row[13][1] ),
    .A1(\second_row[13][1] ),
    .S(_1308_),
    .X(_1311_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1311_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(\first_row[13][0] ),
    .A1(\second_row[13][0] ),
    .S(_1308_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1312_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(\first_row[12][7] ),
    .A1(\second_row[12][7] ),
    .S(_1308_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1313_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(\first_row[12][6] ),
    .A1(\second_row[12][6] ),
    .S(_1308_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _3048_ (.A(_1314_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(\first_row[12][5] ),
    .A1(\second_row[12][5] ),
    .S(_1308_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _3050_ (.A(_1315_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(\first_row[12][4] ),
    .A1(\second_row[12][4] ),
    .S(_1308_),
    .X(_1316_));
 sky130_fd_sc_hd__clkbuf_1 _3052_ (.A(_1316_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(\first_row[12][3] ),
    .A1(\second_row[12][3] ),
    .S(_1308_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_1 _3054_ (.A(_1317_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(\first_row[12][2] ),
    .A1(\second_row[12][2] ),
    .S(_1308_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1318_),
    .X(_0869_));
 sky130_fd_sc_hd__buf_4 _3057_ (.A(_1241_),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(\first_row[12][1] ),
    .A1(\second_row[12][1] ),
    .S(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _3059_ (.A(_1320_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(\first_row[12][0] ),
    .A1(\second_row[12][0] ),
    .S(_1319_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _3061_ (.A(_1321_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(\first_row[11][7] ),
    .A1(\second_row[11][7] ),
    .S(_1319_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _3063_ (.A(_1322_),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(\first_row[11][6] ),
    .A1(\second_row[11][6] ),
    .S(_1319_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _3065_ (.A(_1323_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(\first_row[11][5] ),
    .A1(\second_row[11][5] ),
    .S(_1319_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _3067_ (.A(_1324_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(\first_row[11][4] ),
    .A1(\second_row[11][4] ),
    .S(_1319_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1325_),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(\first_row[11][3] ),
    .A1(\second_row[11][3] ),
    .S(_1319_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_1326_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(\first_row[11][2] ),
    .A1(\second_row[11][2] ),
    .S(_1319_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1327_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(\first_row[11][1] ),
    .A1(\second_row[11][1] ),
    .S(_1319_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1328_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(\first_row[11][0] ),
    .A1(\second_row[11][0] ),
    .S(_1319_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1329_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_4 _3078_ (.A(_1241_),
    .X(_1330_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(\first_row[10][7] ),
    .A1(\second_row[10][7] ),
    .S(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1331_),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(\first_row[10][6] ),
    .A1(\second_row[10][6] ),
    .S(_1330_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _3082_ (.A(_1332_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(\first_row[10][5] ),
    .A1(\second_row[10][5] ),
    .S(_1330_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1333_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(\first_row[10][4] ),
    .A1(\second_row[10][4] ),
    .S(_1330_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_1334_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(\first_row[10][3] ),
    .A1(\second_row[10][3] ),
    .S(_1330_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _3088_ (.A(_1335_),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(\first_row[10][2] ),
    .A1(\second_row[10][2] ),
    .S(_1330_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _3090_ (.A(_1336_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(\first_row[10][1] ),
    .A1(\second_row[10][1] ),
    .S(_1330_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _3092_ (.A(_1337_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(\first_row[10][0] ),
    .A1(\second_row[10][0] ),
    .S(_1330_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1338_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(\first_row[9][7] ),
    .A1(\second_row[9][7] ),
    .S(_1330_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_1339_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(\first_row[9][6] ),
    .A1(\second_row[9][6] ),
    .S(_1330_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1340_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_4 _3099_ (.A(_1241_),
    .X(_1341_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(\first_row[9][5] ),
    .A1(\second_row[9][5] ),
    .S(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _3101_ (.A(_1342_),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(\first_row[9][4] ),
    .A1(\second_row[9][4] ),
    .S(_1341_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _3103_ (.A(_1343_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(\first_row[9][3] ),
    .A1(\second_row[9][3] ),
    .S(_1341_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _3105_ (.A(_1344_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(\first_row[9][2] ),
    .A1(\second_row[9][2] ),
    .S(_1341_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _3107_ (.A(_1345_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(\first_row[9][1] ),
    .A1(\second_row[9][1] ),
    .S(_1341_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _3109_ (.A(_1346_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(\first_row[9][0] ),
    .A1(\second_row[9][0] ),
    .S(_1341_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1347_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(\first_row[8][7] ),
    .A1(\second_row[8][7] ),
    .S(_1341_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1348_),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(\first_row[8][6] ),
    .A1(\second_row[8][6] ),
    .S(_1341_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _3115_ (.A(_1349_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(\first_row[8][5] ),
    .A1(\second_row[8][5] ),
    .S(_1341_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _3117_ (.A(_1350_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(\first_row[8][4] ),
    .A1(\second_row[8][4] ),
    .S(_1341_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _3119_ (.A(_1351_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_4 _3120_ (.A(_1081_),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(\first_row[8][3] ),
    .A1(\second_row[8][3] ),
    .S(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_1353_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(\first_row[8][2] ),
    .A1(\second_row[8][2] ),
    .S(_1352_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _3124_ (.A(_1354_),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(\first_row[8][1] ),
    .A1(\second_row[8][1] ),
    .S(_1352_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1355_),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(\first_row[8][0] ),
    .A1(\second_row[8][0] ),
    .S(_1352_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _3128_ (.A(_1356_),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(\first_row[7][7] ),
    .A1(\second_row[7][7] ),
    .S(_1352_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _3130_ (.A(_1357_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(\first_row[7][6] ),
    .A1(\second_row[7][6] ),
    .S(_1352_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _3132_ (.A(_1358_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(\first_row[7][5] ),
    .A1(\second_row[7][5] ),
    .S(_1352_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _3134_ (.A(_1359_),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(\first_row[7][4] ),
    .A1(\second_row[7][4] ),
    .S(_1352_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _3136_ (.A(_1360_),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(\first_row[7][3] ),
    .A1(\second_row[7][3] ),
    .S(_1352_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _3138_ (.A(_1361_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(\first_row[7][2] ),
    .A1(\second_row[7][2] ),
    .S(_1352_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1362_),
    .X(_0829_));
 sky130_fd_sc_hd__buf_4 _3141_ (.A(_1081_),
    .X(_1363_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(\first_row[7][1] ),
    .A1(\second_row[7][1] ),
    .S(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _3143_ (.A(_1364_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(\first_row[7][0] ),
    .A1(\second_row[7][0] ),
    .S(_1363_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1365_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(\first_row[6][7] ),
    .A1(\second_row[6][7] ),
    .S(_1363_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _3147_ (.A(_1366_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\first_row[6][6] ),
    .A1(\second_row[6][6] ),
    .S(_1363_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1367_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(\first_row[6][5] ),
    .A1(\second_row[6][5] ),
    .S(_1363_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1368_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(\first_row[6][4] ),
    .A1(\second_row[6][4] ),
    .S(_1363_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _3153_ (.A(_1369_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(\first_row[6][3] ),
    .A1(\second_row[6][3] ),
    .S(_1363_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _3155_ (.A(_1370_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(\first_row[6][2] ),
    .A1(\second_row[6][2] ),
    .S(_1363_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _3157_ (.A(_1371_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(\first_row[6][1] ),
    .A1(\second_row[6][1] ),
    .S(_1363_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1372_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(\first_row[6][0] ),
    .A1(\second_row[6][0] ),
    .S(_1363_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _3161_ (.A(_1373_),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _3162_ (.A(_1081_),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(\first_row[5][7] ),
    .A1(\second_row[5][7] ),
    .S(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3164_ (.A(_1375_),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(\first_row[5][6] ),
    .A1(\second_row[5][6] ),
    .S(_1374_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _3166_ (.A(_1376_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\first_row[5][5] ),
    .A1(\second_row[5][5] ),
    .S(_1374_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1377_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\first_row[5][4] ),
    .A1(\second_row[5][4] ),
    .S(_1374_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1378_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(\first_row[5][3] ),
    .A1(\second_row[5][3] ),
    .S(_1374_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1379_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(\first_row[5][2] ),
    .A1(\second_row[5][2] ),
    .S(_1374_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1380_),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\first_row[5][1] ),
    .A1(\second_row[5][1] ),
    .S(_1374_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _3176_ (.A(_1381_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(\first_row[5][0] ),
    .A1(\second_row[5][0] ),
    .S(_1374_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_1382_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(\first_row[4][7] ),
    .A1(\second_row[4][7] ),
    .S(_1374_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _3180_ (.A(_1383_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(\first_row[4][6] ),
    .A1(\second_row[4][6] ),
    .S(_1374_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3182_ (.A(_1384_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_4 _3183_ (.A(_1081_),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(\first_row[4][5] ),
    .A1(\second_row[4][5] ),
    .S(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _3185_ (.A(_1386_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(\first_row[4][4] ),
    .A1(\second_row[4][4] ),
    .S(_1385_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1387_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(\first_row[4][3] ),
    .A1(\second_row[4][3] ),
    .S(_1385_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1388_),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\first_row[4][2] ),
    .A1(\second_row[4][2] ),
    .S(_1385_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1389_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(\first_row[4][1] ),
    .A1(\second_row[4][1] ),
    .S(_1385_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1390_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(\first_row[4][0] ),
    .A1(\second_row[4][0] ),
    .S(_1385_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _3195_ (.A(_1391_),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(\first_row[3][7] ),
    .A1(\second_row[3][7] ),
    .S(_1385_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_1392_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(\first_row[3][6] ),
    .A1(\second_row[3][6] ),
    .S(_1385_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3199_ (.A(_1393_),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(\first_row[3][5] ),
    .A1(\second_row[3][5] ),
    .S(_1385_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3201_ (.A(_1394_),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(\first_row[3][4] ),
    .A1(\second_row[3][4] ),
    .S(_1385_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1395_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_4 _3204_ (.A(_1081_),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(\first_row[3][3] ),
    .A1(\second_row[3][3] ),
    .S(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _3206_ (.A(_1397_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(\first_row[3][2] ),
    .A1(\second_row[3][2] ),
    .S(_1396_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _3208_ (.A(_1398_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(\first_row[3][1] ),
    .A1(\second_row[3][1] ),
    .S(_1396_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1399_),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\first_row[3][0] ),
    .A1(\second_row[3][0] ),
    .S(_1396_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3212_ (.A(_1400_),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\first_row[2][7] ),
    .A1(\second_row[2][7] ),
    .S(_1396_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1401_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\first_row[2][6] ),
    .A1(\second_row[2][6] ),
    .S(_1396_),
    .X(_1402_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1402_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\first_row[2][5] ),
    .A1(\second_row[2][5] ),
    .S(_1396_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _3218_ (.A(_1403_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\first_row[2][4] ),
    .A1(\second_row[2][4] ),
    .S(_1396_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _3220_ (.A(_1404_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\first_row[2][3] ),
    .A1(\second_row[2][3] ),
    .S(_1396_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3222_ (.A(_1405_),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\first_row[2][2] ),
    .A1(\second_row[2][2] ),
    .S(_1396_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1406_),
    .X(_0789_));
 sky130_fd_sc_hd__buf_4 _3225_ (.A(_1081_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(\first_row[2][1] ),
    .A1(\second_row[2][1] ),
    .S(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3227_ (.A(_1408_),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\first_row[2][0] ),
    .A1(\second_row[2][0] ),
    .S(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _3229_ (.A(_1409_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\first_row[1][7] ),
    .A1(\second_row[1][7] ),
    .S(_1407_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _3231_ (.A(_1410_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(\first_row[1][6] ),
    .A1(\second_row[1][6] ),
    .S(_1407_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _3233_ (.A(_1411_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(\first_row[1][5] ),
    .A1(\second_row[1][5] ),
    .S(_1407_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_1412_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(\first_row[1][4] ),
    .A1(\second_row[1][4] ),
    .S(_1407_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3237_ (.A(_1413_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(\first_row[1][3] ),
    .A1(\second_row[1][3] ),
    .S(_1407_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3239_ (.A(_1414_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(\first_row[1][2] ),
    .A1(\second_row[1][2] ),
    .S(_1407_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_1415_),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(\first_row[1][1] ),
    .A1(\second_row[1][1] ),
    .S(_1407_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _3243_ (.A(_1416_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(\first_row[1][0] ),
    .A1(\second_row[1][0] ),
    .S(_1407_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _3245_ (.A(_1417_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(\first_row[0][7] ),
    .A1(\second_row[0][7] ),
    .S(_1082_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_1418_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(\first_row[0][6] ),
    .A1(\second_row[0][6] ),
    .S(_1082_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3249_ (.A(_1419_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(\first_row[0][5] ),
    .A1(\second_row[0][5] ),
    .S(_1082_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3251_ (.A(_1420_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(\first_row[0][4] ),
    .A1(\second_row[0][4] ),
    .S(_1082_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1421_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(\first_row[0][3] ),
    .A1(\second_row[0][3] ),
    .S(_1082_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1422_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\first_row[0][2] ),
    .A1(\second_row[0][2] ),
    .S(_1082_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_1423_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(\first_row[0][1] ),
    .A1(\second_row[0][1] ),
    .S(_1082_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1424_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(\first_row[0][0] ),
    .A1(\second_row[0][0] ),
    .S(_1082_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1425_),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _3262_ (.A(_1067_),
    .B(_1098_),
    .X(_1426_));
 sky130_fd_sc_hd__buf_2 _3263_ (.A(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__or3_1 _3264_ (.A(_1094_),
    .B(_1078_),
    .C(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_4 _3265_ (.A(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(_1092_),
    .A1(\first_row[17][7] ),
    .S(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3267_ (.A(_1430_),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(_1103_),
    .A1(\first_row[17][6] ),
    .S(_1429_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3269_ (.A(_1431_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(_1105_),
    .A1(\first_row[17][5] ),
    .S(_1429_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_1432_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(_1107_),
    .A1(\first_row[17][4] ),
    .S(_1429_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1433_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(_1109_),
    .A1(\first_row[17][3] ),
    .S(_1429_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3275_ (.A(_1434_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(_1111_),
    .A1(\first_row[17][2] ),
    .S(_1429_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3277_ (.A(_1435_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(_1113_),
    .A1(\first_row[17][1] ),
    .S(_1429_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1436_),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(_1115_),
    .A1(\first_row[17][0] ),
    .S(_1429_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _3281_ (.A(_1437_),
    .X(_0763_));
 sky130_fd_sc_hd__and4_1 _3282_ (.A(\col_input[4] ),
    .B(_1093_),
    .C(_1095_),
    .D(_1099_),
    .X(_1438_));
 sky130_fd_sc_hd__buf_2 _3283_ (.A(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\first_row[16][7] ),
    .A1(net8),
    .S(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3285_ (.A(_1440_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(\first_row[16][6] ),
    .A1(net7),
    .S(_1439_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_1 _3287_ (.A(_1441_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\first_row[16][5] ),
    .A1(net6),
    .S(_1439_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1442_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\first_row[16][4] ),
    .A1(net5),
    .S(_1439_),
    .X(_1443_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1443_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\first_row[16][3] ),
    .A1(net4),
    .S(_1439_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1444_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(\first_row[16][2] ),
    .A1(net3),
    .S(_1439_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3295_ (.A(_1445_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(\first_row[16][1] ),
    .A1(net2),
    .S(_1439_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(_1446_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(\first_row[16][0] ),
    .A1(net1),
    .S(_1439_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(_1447_),
    .X(_0755_));
 sky130_fd_sc_hd__inv_2 _3300_ (.A(\col_input[1] ),
    .Y(_1448_));
 sky130_fd_sc_hd__or4b_2 _3301_ (.A(_1067_),
    .B(_1448_),
    .C(_1098_),
    .D_N(\col_input[0] ),
    .X(_1449_));
 sky130_fd_sc_hd__nand2_1 _3302_ (.A(_1077_),
    .B(\col_input[2] ),
    .Y(_1450_));
 sky130_fd_sc_hd__nor2_1 _3303_ (.A(_1449_),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_4 _3304_ (.A(_1094_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(_1092_),
    .A1(\first_row[15][7] ),
    .S(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _3306_ (.A(_1453_),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_1103_),
    .A1(\first_row[15][6] ),
    .S(_1452_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(_1454_),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(_1105_),
    .A1(\first_row[15][5] ),
    .S(_1452_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1455_),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(_1107_),
    .A1(\first_row[15][4] ),
    .S(_1452_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _3312_ (.A(_1456_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(_1109_),
    .A1(\first_row[15][3] ),
    .S(_1452_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3314_ (.A(_1457_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(_1111_),
    .A1(\first_row[15][2] ),
    .S(_1452_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1458_),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(_1113_),
    .A1(\first_row[15][1] ),
    .S(_1452_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3318_ (.A(_1459_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(_1115_),
    .A1(\first_row[15][0] ),
    .S(_1452_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _3320_ (.A(_1460_),
    .X(_0747_));
 sky130_fd_sc_hd__or4_1 _3321_ (.A(\col_input[4] ),
    .B(_1448_),
    .C(\col_input[0] ),
    .D(_1427_),
    .X(_1461_));
 sky130_fd_sc_hd__or2_1 _3322_ (.A(_1450_),
    .B(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_4 _3323_ (.A(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(_1092_),
    .A1(\first_row[14][7] ),
    .S(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1464_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(_1103_),
    .A1(\first_row[14][6] ),
    .S(_1463_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3327_ (.A(_1465_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(_1105_),
    .A1(\first_row[14][5] ),
    .S(_1463_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1466_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(_1107_),
    .A1(\first_row[14][4] ),
    .S(_1463_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3331_ (.A(_1467_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(_1109_),
    .A1(\first_row[14][3] ),
    .S(_1463_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3333_ (.A(_1468_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(_1111_),
    .A1(\first_row[14][2] ),
    .S(_1463_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3335_ (.A(_1469_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _3336_ (.A0(_1113_),
    .A1(\first_row[14][1] ),
    .S(_1463_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _3337_ (.A(_1470_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(_1115_),
    .A1(\first_row[14][0] ),
    .S(_1463_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3339_ (.A(_1471_),
    .X(_0739_));
 sky130_fd_sc_hd__or4b_1 _3340_ (.A(\col_input[4] ),
    .B(_1427_),
    .C(\col_input[1] ),
    .D_N(\col_input[0] ),
    .X(_1472_));
 sky130_fd_sc_hd__or2_1 _3341_ (.A(_1450_),
    .B(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_4 _3342_ (.A(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(_1092_),
    .A1(\first_row[13][7] ),
    .S(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3344_ (.A(_1475_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(_1103_),
    .A1(\first_row[13][6] ),
    .S(_1474_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3346_ (.A(_1476_),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(_1105_),
    .A1(\first_row[13][5] ),
    .S(_1474_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3348_ (.A(_1477_),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(_1107_),
    .A1(\first_row[13][4] ),
    .S(_1474_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3350_ (.A(_1478_),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(_1109_),
    .A1(\first_row[13][3] ),
    .S(_1474_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3352_ (.A(_1479_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(_1111_),
    .A1(\first_row[13][2] ),
    .S(_1474_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3354_ (.A(_1480_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(_1113_),
    .A1(\first_row[13][1] ),
    .S(_1474_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3356_ (.A(_1481_),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(_1115_),
    .A1(\first_row[13][0] ),
    .S(_1474_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3358_ (.A(_1482_),
    .X(_0731_));
 sky130_fd_sc_hd__and2_1 _3359_ (.A(_1077_),
    .B(\col_input[2] ),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_4 _3360_ (.A(_1100_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(_1092_),
    .A1(\first_row[12][7] ),
    .S(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(_1485_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(_1103_),
    .A1(\first_row[12][6] ),
    .S(_1484_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3364_ (.A(_1486_),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(_1105_),
    .A1(\first_row[12][5] ),
    .S(_1484_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(_1487_),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(_1107_),
    .A1(\first_row[12][4] ),
    .S(_1484_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3368_ (.A(_1488_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(_1109_),
    .A1(\first_row[12][3] ),
    .S(_1484_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _3370_ (.A(_1489_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(_1111_),
    .A1(\first_row[12][2] ),
    .S(_1484_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1490_),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(_1113_),
    .A1(\first_row[12][1] ),
    .S(_1484_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1491_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(_1115_),
    .A1(\first_row[12][0] ),
    .S(_1484_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_1 _3376_ (.A(_1492_),
    .X(_0723_));
 sky130_fd_sc_hd__nor2_2 _3377_ (.A(\col_input[4] ),
    .B(_1449_),
    .Y(_1493_));
 sky130_fd_sc_hd__inv_2 _3378_ (.A(\col_input[2] ),
    .Y(_1494_));
 sky130_fd_sc_hd__and2_4 _3379_ (.A(_1077_),
    .B(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nand2_4 _3380_ (.A(_1493_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(_1092_),
    .A1(\first_row[11][7] ),
    .S(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _3382_ (.A(_1497_),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(_1103_),
    .A1(\first_row[11][6] ),
    .S(_1496_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3384_ (.A(_1498_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(_1105_),
    .A1(\first_row[11][5] ),
    .S(_1496_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3386_ (.A(_1499_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(_1107_),
    .A1(\first_row[11][4] ),
    .S(_1496_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3388_ (.A(_1500_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(_1109_),
    .A1(\first_row[11][3] ),
    .S(_1496_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3390_ (.A(_1501_),
    .X(_0718_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(_1111_),
    .A1(\first_row[11][2] ),
    .S(_1496_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3392_ (.A(_1502_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(_1113_),
    .A1(\first_row[11][1] ),
    .S(_1496_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3394_ (.A(_1503_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(_1115_),
    .A1(\first_row[11][0] ),
    .S(_1496_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3396_ (.A(_1504_),
    .X(_0715_));
 sky130_fd_sc_hd__nand2b_4 _3397_ (.A_N(_1461_),
    .B(_1495_),
    .Y(_1505_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(_1092_),
    .A1(\first_row[10][7] ),
    .S(_1505_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3399_ (.A(_1506_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(_1103_),
    .A1(\first_row[10][6] ),
    .S(_1505_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3401_ (.A(_1507_),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(_1105_),
    .A1(\first_row[10][5] ),
    .S(_1505_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _3403_ (.A(_1508_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(_1107_),
    .A1(\first_row[10][4] ),
    .S(_1505_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _3405_ (.A(_1509_),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(_1109_),
    .A1(\first_row[10][3] ),
    .S(_1505_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3407_ (.A(_1510_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(_1111_),
    .A1(\first_row[10][2] ),
    .S(_1505_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3409_ (.A(_1511_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(_1113_),
    .A1(\first_row[10][1] ),
    .S(_1505_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3411_ (.A(_1512_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(_1115_),
    .A1(\first_row[10][0] ),
    .S(_1505_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3413_ (.A(_1513_),
    .X(_0707_));
 sky130_fd_sc_hd__nand2b_4 _3414_ (.A_N(_1472_),
    .B(_1495_),
    .Y(_1514_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(_1092_),
    .A1(\first_row[9][7] ),
    .S(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3416_ (.A(_1515_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(_1103_),
    .A1(\first_row[9][6] ),
    .S(_1514_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3418_ (.A(_1516_),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(_1105_),
    .A1(\first_row[9][5] ),
    .S(_1514_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3420_ (.A(_1517_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(_1107_),
    .A1(\first_row[9][4] ),
    .S(_1514_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3422_ (.A(_1518_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(_1109_),
    .A1(\first_row[9][3] ),
    .S(_1514_),
    .X(_1519_));
 sky130_fd_sc_hd__clkbuf_1 _3424_ (.A(_1519_),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(_1111_),
    .A1(\first_row[9][2] ),
    .S(_1514_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3426_ (.A(_1520_),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(_1113_),
    .A1(\first_row[9][1] ),
    .S(_1514_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3428_ (.A(_1521_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(_1115_),
    .A1(\first_row[9][0] ),
    .S(_1514_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3430_ (.A(_1522_),
    .X(_0699_));
 sky130_fd_sc_hd__nand2_4 _3431_ (.A(_1100_),
    .B(_1495_),
    .Y(_1523_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(_1092_),
    .A1(\first_row[8][7] ),
    .S(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3433_ (.A(_1524_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(_1103_),
    .A1(\first_row[8][6] ),
    .S(_1523_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _3435_ (.A(_1525_),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(_1105_),
    .A1(\first_row[8][5] ),
    .S(_1523_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3437_ (.A(_1526_),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(_1107_),
    .A1(\first_row[8][4] ),
    .S(_1523_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3439_ (.A(_1527_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(_1109_),
    .A1(\first_row[8][3] ),
    .S(_1523_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3441_ (.A(_1528_),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(_1111_),
    .A1(\first_row[8][2] ),
    .S(_1523_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3443_ (.A(_1529_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(_1113_),
    .A1(\first_row[8][1] ),
    .S(_1523_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3445_ (.A(_1530_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(_1115_),
    .A1(\first_row[8][0] ),
    .S(_1523_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3447_ (.A(_1531_),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_2 _3448_ (.A(_1077_),
    .B(_1494_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_4 _3449_ (.A(_1493_),
    .B(_1532_),
    .Y(_1533_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(net8),
    .A1(\first_row[7][7] ),
    .S(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3451_ (.A(_1534_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(net7),
    .A1(\first_row[7][6] ),
    .S(_1533_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3453_ (.A(_1535_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(net6),
    .A1(\first_row[7][5] ),
    .S(_1533_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3455_ (.A(_1536_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(net5),
    .A1(\first_row[7][4] ),
    .S(_1533_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3457_ (.A(_1537_),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(net4),
    .A1(\first_row[7][3] ),
    .S(_1533_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3459_ (.A(_1538_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(net3),
    .A1(\first_row[7][2] ),
    .S(_1533_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3461_ (.A(_1539_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(net2),
    .A1(\first_row[7][1] ),
    .S(_1533_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3463_ (.A(_1540_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(net1),
    .A1(\first_row[7][0] ),
    .S(_1533_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1541_),
    .X(_0683_));
 sky130_fd_sc_hd__or3_2 _3466_ (.A(_1077_),
    .B(_1494_),
    .C(_1461_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_4 _3467_ (.A(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(net8),
    .A1(\first_row[6][7] ),
    .S(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3469_ (.A(_1544_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(net7),
    .A1(\first_row[6][6] ),
    .S(_1543_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3471_ (.A(_1545_),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(net6),
    .A1(\first_row[6][5] ),
    .S(_1543_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_1 _3473_ (.A(_1546_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(net5),
    .A1(\first_row[6][4] ),
    .S(_1543_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3475_ (.A(_1547_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(net4),
    .A1(\first_row[6][3] ),
    .S(_1543_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _3477_ (.A(_1548_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(net3),
    .A1(\first_row[6][2] ),
    .S(_1543_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3479_ (.A(_1549_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(net2),
    .A1(\first_row[6][1] ),
    .S(_1543_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _3481_ (.A(_1550_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(net1),
    .A1(\first_row[6][0] ),
    .S(_1543_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3483_ (.A(_1551_),
    .X(_0675_));
 sky130_fd_sc_hd__or3_2 _3484_ (.A(_1077_),
    .B(_1494_),
    .C(_1472_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_4 _3485_ (.A(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(net8),
    .A1(\first_row[5][7] ),
    .S(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _3487_ (.A(_1554_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(net7),
    .A1(\first_row[5][6] ),
    .S(_1553_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3489_ (.A(_1555_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(net6),
    .A1(\first_row[5][5] ),
    .S(_1553_),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _3491_ (.A(_1556_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(net5),
    .A1(\first_row[5][4] ),
    .S(_1553_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3493_ (.A(_1557_),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(net4),
    .A1(\first_row[5][3] ),
    .S(_1553_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3495_ (.A(_1558_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(net3),
    .A1(\first_row[5][2] ),
    .S(_1553_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3497_ (.A(_1559_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(net2),
    .A1(\first_row[5][1] ),
    .S(_1553_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1560_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(net1),
    .A1(\first_row[5][0] ),
    .S(_1553_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(_1561_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_8 _3502_ (.A(_1100_),
    .B(_1532_),
    .Y(_1562_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(net8),
    .A1(\first_row[4][7] ),
    .S(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _3504_ (.A(_1563_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(net7),
    .A1(\first_row[4][6] ),
    .S(_1562_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3506_ (.A(_1564_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(net6),
    .A1(\first_row[4][5] ),
    .S(_1562_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(_1565_),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(net5),
    .A1(\first_row[4][4] ),
    .S(_1562_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_1566_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(net4),
    .A1(\first_row[4][3] ),
    .S(_1562_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3512_ (.A(_1567_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(net3),
    .A1(\first_row[4][2] ),
    .S(_1562_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3514_ (.A(_1568_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(net2),
    .A1(\first_row[4][1] ),
    .S(_1562_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3516_ (.A(_1569_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(net1),
    .A1(\first_row[4][0] ),
    .S(_1562_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3518_ (.A(_1570_),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_4 _3519_ (.A(_1093_),
    .B(_1493_),
    .Y(_1571_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(net8),
    .A1(\first_row[3][7] ),
    .S(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _3521_ (.A(_1572_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(net7),
    .A1(\first_row[3][6] ),
    .S(_1571_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3523_ (.A(_1573_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(net6),
    .A1(\first_row[3][5] ),
    .S(_1571_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3525_ (.A(_1574_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(net5),
    .A1(\first_row[3][4] ),
    .S(_1571_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3527_ (.A(_1575_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(net4),
    .A1(\first_row[3][3] ),
    .S(_1571_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3529_ (.A(_1576_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(net3),
    .A1(\first_row[3][2] ),
    .S(_1571_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3531_ (.A(_1577_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(net2),
    .A1(\first_row[3][1] ),
    .S(_1571_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3533_ (.A(_1578_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(net1),
    .A1(\first_row[3][0] ),
    .S(_1571_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3535_ (.A(_1579_),
    .X(_0651_));
 sky130_fd_sc_hd__or3_1 _3536_ (.A(_1077_),
    .B(\col_input[2] ),
    .C(_1461_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_4 _3537_ (.A(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(net8),
    .A1(\first_row[2][7] ),
    .S(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3539_ (.A(_1582_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _3540_ (.A0(net7),
    .A1(\first_row[2][6] ),
    .S(_1581_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3541_ (.A(_1583_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(net6),
    .A1(\first_row[2][5] ),
    .S(_1581_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3543_ (.A(_1584_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(net5),
    .A1(\first_row[2][4] ),
    .S(_1581_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3545_ (.A(_1585_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(net4),
    .A1(\first_row[2][3] ),
    .S(_1581_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3547_ (.A(_1586_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(net3),
    .A1(\first_row[2][2] ),
    .S(_1581_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3549_ (.A(_1587_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(net2),
    .A1(\first_row[2][1] ),
    .S(_1581_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1588_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(net1),
    .A1(\first_row[2][0] ),
    .S(_1581_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1589_),
    .X(_0643_));
 sky130_fd_sc_hd__or3_1 _3554_ (.A(_1077_),
    .B(\col_input[2] ),
    .C(_1472_),
    .X(_1590_));
 sky130_fd_sc_hd__buf_4 _3555_ (.A(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(net8),
    .A1(\first_row[1][7] ),
    .S(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3557_ (.A(_1592_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(net7),
    .A1(\first_row[1][6] ),
    .S(_1591_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3559_ (.A(_1593_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(net6),
    .A1(\first_row[1][5] ),
    .S(_1591_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3561_ (.A(_1594_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(net5),
    .A1(\first_row[1][4] ),
    .S(_1591_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3563_ (.A(_1595_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(net4),
    .A1(\first_row[1][3] ),
    .S(_1591_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3565_ (.A(_1596_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(net3),
    .A1(\first_row[1][2] ),
    .S(_1591_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3567_ (.A(_1597_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(net2),
    .A1(\first_row[1][1] ),
    .S(_1591_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3569_ (.A(_1598_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(net1),
    .A1(\first_row[1][0] ),
    .S(_1591_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3571_ (.A(_1599_),
    .X(_0635_));
 sky130_fd_sc_hd__or4_1 _3572_ (.A(\k[26] ),
    .B(\k[25] ),
    .C(\k[24] ),
    .D(\k[23] ),
    .X(_1600_));
 sky130_fd_sc_hd__or4_1 _3573_ (.A(\k[18] ),
    .B(\k[17] ),
    .C(\k[16] ),
    .D(\k[15] ),
    .X(_1601_));
 sky130_fd_sc_hd__or4_1 _3574_ (.A(\k[22] ),
    .B(\k[21] ),
    .C(\k[20] ),
    .D(\k[19] ),
    .X(_1602_));
 sky130_fd_sc_hd__or4_1 _3575_ (.A(\k[14] ),
    .B(\k[13] ),
    .C(\k[12] ),
    .D(\k[11] ),
    .X(_1603_));
 sky130_fd_sc_hd__or4_1 _3576_ (.A(\k[10] ),
    .B(\k[9] ),
    .C(\k[8] ),
    .D(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__or4_1 _3577_ (.A(\k[30] ),
    .B(\k[29] ),
    .C(\k[28] ),
    .D(\k[27] ),
    .X(_1605_));
 sky130_fd_sc_hd__or4_1 _3578_ (.A(_1601_),
    .B(_1602_),
    .C(_1604_),
    .D(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__o21bai_1 _3579_ (.A1(_1600_),
    .A2(_1606_),
    .B1_N(\k[31] ),
    .Y(_1607_));
 sky130_fd_sc_hd__or3_1 _3580_ (.A(\valid_counter[6] ),
    .B(\valid_counter[5] ),
    .C(\valid_counter[4] ),
    .X(_1608_));
 sky130_fd_sc_hd__or4_1 _3581_ (.A(\valid_counter[10] ),
    .B(\valid_counter[9] ),
    .C(\valid_counter[8] ),
    .D(\valid_counter[7] ),
    .X(_1609_));
 sky130_fd_sc_hd__or4_1 _3582_ (.A(\valid_counter[14] ),
    .B(\valid_counter[13] ),
    .C(\valid_counter[12] ),
    .D(\valid_counter[11] ),
    .X(_1610_));
 sky130_fd_sc_hd__or4_1 _3583_ (.A(\valid_counter[26] ),
    .B(\valid_counter[25] ),
    .C(\valid_counter[24] ),
    .D(\valid_counter[23] ),
    .X(_1611_));
 sky130_fd_sc_hd__or4_1 _3584_ (.A(\valid_counter[30] ),
    .B(\valid_counter[29] ),
    .C(\valid_counter[28] ),
    .D(\valid_counter[27] ),
    .X(_1612_));
 sky130_fd_sc_hd__or4_1 _3585_ (.A(\valid_counter[18] ),
    .B(\valid_counter[17] ),
    .C(\valid_counter[16] ),
    .D(\valid_counter[15] ),
    .X(_1613_));
 sky130_fd_sc_hd__or4_1 _3586_ (.A(\valid_counter[22] ),
    .B(\valid_counter[21] ),
    .C(\valid_counter[20] ),
    .D(\valid_counter[19] ),
    .X(_1614_));
 sky130_fd_sc_hd__or4_1 _3587_ (.A(_1611_),
    .B(_1612_),
    .C(_1613_),
    .D(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__or4_1 _3588_ (.A(_1608_),
    .B(_1609_),
    .C(_1610_),
    .D(_1615_),
    .X(_1616_));
 sky130_fd_sc_hd__and3b_1 _3589_ (.A_N(\valid_counter[31] ),
    .B(_1607_),
    .C(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__or4_1 _3590_ (.A(\k[3] ),
    .B(\k[2] ),
    .C(\k[1] ),
    .D(\k[0] ),
    .X(_1618_));
 sky130_fd_sc_hd__or4_1 _3591_ (.A(\k[7] ),
    .B(\k[6] ),
    .C(\k[5] ),
    .D(\k[4] ),
    .X(_1619_));
 sky130_fd_sc_hd__nor2_1 _3592_ (.A(_1618_),
    .B(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hd__o211ai_1 _3593_ (.A1(\k[31] ),
    .A2(_1620_),
    .B1(_1607_),
    .C1(_1067_),
    .Y(_1621_));
 sky130_fd_sc_hd__o2111a_1 _3594_ (.A1(_1067_),
    .A2(_1617_),
    .B1(_1621_),
    .C1(\k[1] ),
    .D1(\k[0] ),
    .X(_1622_));
 sky130_fd_sc_hd__and4_1 _3595_ (.A(\k[4] ),
    .B(\k[3] ),
    .C(\k[2] ),
    .D(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__and4_1 _3596_ (.A(\k[7] ),
    .B(\k[6] ),
    .C(\k[5] ),
    .D(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and4_1 _3597_ (.A(\k[10] ),
    .B(\k[9] ),
    .C(\k[8] ),
    .D(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__and4_1 _3598_ (.A(\k[13] ),
    .B(\k[12] ),
    .C(\k[11] ),
    .D(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__and4_1 _3599_ (.A(\k[16] ),
    .B(\k[15] ),
    .C(\k[14] ),
    .D(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__and4_1 _3600_ (.A(\k[19] ),
    .B(\k[18] ),
    .C(\k[17] ),
    .D(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__and3_1 _3601_ (.A(\k[21] ),
    .B(\k[20] ),
    .C(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__and2_1 _3602_ (.A(\k[22] ),
    .B(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__and3_1 _3603_ (.A(\k[24] ),
    .B(\k[23] ),
    .C(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__and2_1 _3604_ (.A(\k[25] ),
    .B(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__and3_1 _3605_ (.A(\k[27] ),
    .B(\k[26] ),
    .C(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__and2_1 _3606_ (.A(\k[28] ),
    .B(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__and3_1 _3607_ (.A(\k[30] ),
    .B(\k[29] ),
    .C(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__xor2_1 _3608_ (.A(\k[31] ),
    .B(_1635_),
    .X(_0634_));
 sky130_fd_sc_hd__a21oi_1 _3609_ (.A1(\k[29] ),
    .A2(_1634_),
    .B1(\k[30] ),
    .Y(_1636_));
 sky130_fd_sc_hd__nor2_1 _3610_ (.A(_1635_),
    .B(_1636_),
    .Y(_0633_));
 sky130_fd_sc_hd__xor2_1 _3611_ (.A(\k[29] ),
    .B(_1634_),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_1 _3612_ (.A(\k[28] ),
    .B(_1633_),
    .Y(_1637_));
 sky130_fd_sc_hd__nor2_1 _3613_ (.A(_1634_),
    .B(_1637_),
    .Y(_0631_));
 sky130_fd_sc_hd__a31o_1 _3614_ (.A1(\k[26] ),
    .A2(\k[25] ),
    .A3(_1631_),
    .B1(\k[27] ),
    .X(_1638_));
 sky130_fd_sc_hd__and2b_1 _3615_ (.A_N(_1633_),
    .B(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _3616_ (.A(_1639_),
    .X(_0630_));
 sky130_fd_sc_hd__xor2_1 _3617_ (.A(\k[26] ),
    .B(_1632_),
    .X(_0629_));
 sky130_fd_sc_hd__nor2_1 _3618_ (.A(\k[25] ),
    .B(_1631_),
    .Y(_1640_));
 sky130_fd_sc_hd__nor2_1 _3619_ (.A(_1632_),
    .B(_1640_),
    .Y(_0628_));
 sky130_fd_sc_hd__a21oi_1 _3620_ (.A1(\k[23] ),
    .A2(_1630_),
    .B1(\k[24] ),
    .Y(_1641_));
 sky130_fd_sc_hd__nor2_1 _3621_ (.A(_1631_),
    .B(_1641_),
    .Y(_0627_));
 sky130_fd_sc_hd__xor2_1 _3622_ (.A(\k[23] ),
    .B(_1630_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _3623_ (.A(\k[22] ),
    .B(_1629_),
    .Y(_1642_));
 sky130_fd_sc_hd__nor2_1 _3624_ (.A(_1630_),
    .B(_1642_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_1 _3625_ (.A1(\k[20] ),
    .A2(_1628_),
    .B1(\k[21] ),
    .Y(_1643_));
 sky130_fd_sc_hd__nor2_1 _3626_ (.A(_1629_),
    .B(_1643_),
    .Y(_0624_));
 sky130_fd_sc_hd__xor2_1 _3627_ (.A(\k[20] ),
    .B(_1628_),
    .X(_0623_));
 sky130_fd_sc_hd__a31o_1 _3628_ (.A1(\k[18] ),
    .A2(\k[17] ),
    .A3(_1627_),
    .B1(\k[19] ),
    .X(_1644_));
 sky130_fd_sc_hd__and2b_1 _3629_ (.A_N(_1628_),
    .B(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3630_ (.A(_1645_),
    .X(_0622_));
 sky130_fd_sc_hd__nand2_1 _3631_ (.A(\k[17] ),
    .B(_1627_),
    .Y(_1646_));
 sky130_fd_sc_hd__xnor2_1 _3632_ (.A(\k[18] ),
    .B(_1646_),
    .Y(_0621_));
 sky130_fd_sc_hd__xor2_1 _3633_ (.A(\k[17] ),
    .B(_1627_),
    .X(_0620_));
 sky130_fd_sc_hd__a31o_1 _3634_ (.A1(\k[15] ),
    .A2(\k[14] ),
    .A3(_1626_),
    .B1(\k[16] ),
    .X(_1647_));
 sky130_fd_sc_hd__and2b_1 _3635_ (.A_N(_1627_),
    .B(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3636_ (.A(_1648_),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(\k[14] ),
    .B(_1626_),
    .Y(_1649_));
 sky130_fd_sc_hd__xnor2_1 _3638_ (.A(\k[15] ),
    .B(_1649_),
    .Y(_0618_));
 sky130_fd_sc_hd__xor2_1 _3639_ (.A(\k[14] ),
    .B(_1626_),
    .X(_0617_));
 sky130_fd_sc_hd__a31o_1 _3640_ (.A1(\k[12] ),
    .A2(\k[11] ),
    .A3(_1625_),
    .B1(\k[13] ),
    .X(_1650_));
 sky130_fd_sc_hd__and2b_1 _3641_ (.A_N(_1626_),
    .B(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _3642_ (.A(_1651_),
    .X(_0616_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(\k[11] ),
    .B(_1625_),
    .Y(_1652_));
 sky130_fd_sc_hd__xnor2_1 _3644_ (.A(\k[12] ),
    .B(_1652_),
    .Y(_0615_));
 sky130_fd_sc_hd__xor2_1 _3645_ (.A(\k[11] ),
    .B(_1625_),
    .X(_0614_));
 sky130_fd_sc_hd__a31o_1 _3646_ (.A1(\k[9] ),
    .A2(\k[8] ),
    .A3(_1624_),
    .B1(\k[10] ),
    .X(_1653_));
 sky130_fd_sc_hd__and2b_1 _3647_ (.A_N(_1625_),
    .B(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3648_ (.A(_1654_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(\k[8] ),
    .B(_1624_),
    .Y(_1655_));
 sky130_fd_sc_hd__xnor2_1 _3650_ (.A(\k[9] ),
    .B(_1655_),
    .Y(_0612_));
 sky130_fd_sc_hd__xor2_1 _3651_ (.A(\k[8] ),
    .B(_1624_),
    .X(_0611_));
 sky130_fd_sc_hd__a31o_1 _3652_ (.A1(\k[6] ),
    .A2(\k[5] ),
    .A3(_1623_),
    .B1(\k[7] ),
    .X(_1656_));
 sky130_fd_sc_hd__and2b_1 _3653_ (.A_N(_1624_),
    .B(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3654_ (.A(_1657_),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(\k[5] ),
    .B(_1623_),
    .Y(_1658_));
 sky130_fd_sc_hd__xnor2_1 _3656_ (.A(\k[6] ),
    .B(_1658_),
    .Y(_0609_));
 sky130_fd_sc_hd__xor2_1 _3657_ (.A(\k[5] ),
    .B(_1623_),
    .X(_0608_));
 sky130_fd_sc_hd__a31o_1 _3658_ (.A1(\k[3] ),
    .A2(\k[2] ),
    .A3(_1622_),
    .B1(\k[4] ),
    .X(_1659_));
 sky130_fd_sc_hd__and2b_1 _3659_ (.A_N(_1623_),
    .B(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3660_ (.A(_1660_),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _3661_ (.A(\k[2] ),
    .B(_1622_),
    .Y(_1661_));
 sky130_fd_sc_hd__xnor2_1 _3662_ (.A(\k[3] ),
    .B(_1661_),
    .Y(_0606_));
 sky130_fd_sc_hd__or2_1 _3663_ (.A(\k[2] ),
    .B(_1622_),
    .X(_1662_));
 sky130_fd_sc_hd__and2_1 _3664_ (.A(_1661_),
    .B(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3665_ (.A(_1663_),
    .X(_0605_));
 sky130_fd_sc_hd__o21a_1 _3666_ (.A1(_1067_),
    .A2(_1617_),
    .B1(_1621_),
    .X(_1664_));
 sky130_fd_sc_hd__and2_1 _3667_ (.A(\k[0] ),
    .B(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__nor2_1 _3668_ (.A(\k[1] ),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__nor2_1 _3669_ (.A(_1622_),
    .B(_1666_),
    .Y(_0604_));
 sky130_fd_sc_hd__nor2_1 _3670_ (.A(\k[0] ),
    .B(_1664_),
    .Y(_1667_));
 sky130_fd_sc_hd__nor2_1 _3671_ (.A(_1665_),
    .B(_1667_),
    .Y(_0603_));
 sky130_fd_sc_hd__and4_1 _3672_ (.A(net10),
    .B(\valid_counter[2] ),
    .C(\valid_counter[1] ),
    .D(\valid_counter[0] ),
    .X(_1668_));
 sky130_fd_sc_hd__and4_1 _3673_ (.A(\valid_counter[5] ),
    .B(\valid_counter[4] ),
    .C(\valid_counter[3] ),
    .D(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__and3_1 _3674_ (.A(\valid_counter[7] ),
    .B(\valid_counter[6] ),
    .C(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__and2_1 _3675_ (.A(\valid_counter[8] ),
    .B(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__and3_1 _3676_ (.A(\valid_counter[10] ),
    .B(\valid_counter[9] ),
    .C(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__and2_1 _3677_ (.A(\valid_counter[11] ),
    .B(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__and3_1 _3678_ (.A(\valid_counter[13] ),
    .B(\valid_counter[12] ),
    .C(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__and2_1 _3679_ (.A(\valid_counter[14] ),
    .B(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__and3_1 _3680_ (.A(\valid_counter[16] ),
    .B(\valid_counter[15] ),
    .C(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and2_1 _3681_ (.A(\valid_counter[17] ),
    .B(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__and3_1 _3682_ (.A(\valid_counter[19] ),
    .B(\valid_counter[18] ),
    .C(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__and2_1 _3683_ (.A(\valid_counter[20] ),
    .B(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__and3_1 _3684_ (.A(\valid_counter[22] ),
    .B(\valid_counter[21] ),
    .C(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__and2_1 _3685_ (.A(\valid_counter[23] ),
    .B(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__and3_1 _3686_ (.A(\valid_counter[25] ),
    .B(\valid_counter[24] ),
    .C(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__and2_1 _3687_ (.A(\valid_counter[26] ),
    .B(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__and3_1 _3688_ (.A(\valid_counter[28] ),
    .B(\valid_counter[27] ),
    .C(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__and2_1 _3689_ (.A(\valid_counter[29] ),
    .B(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _3690_ (.A(\valid_counter[30] ),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__xnor2_1 _3691_ (.A(\valid_counter[31] ),
    .B(_1686_),
    .Y(_0602_));
 sky130_fd_sc_hd__xor2_1 _3692_ (.A(\valid_counter[30] ),
    .B(_1685_),
    .X(_0601_));
 sky130_fd_sc_hd__nor2_1 _3693_ (.A(\valid_counter[29] ),
    .B(_1684_),
    .Y(_1687_));
 sky130_fd_sc_hd__nor2_1 _3694_ (.A(_1685_),
    .B(_1687_),
    .Y(_0600_));
 sky130_fd_sc_hd__a31o_1 _3695_ (.A1(\valid_counter[27] ),
    .A2(\valid_counter[26] ),
    .A3(_1682_),
    .B1(\valid_counter[28] ),
    .X(_1688_));
 sky130_fd_sc_hd__and2b_1 _3696_ (.A_N(_1684_),
    .B(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3697_ (.A(_1689_),
    .X(_0599_));
 sky130_fd_sc_hd__xor2_1 _3698_ (.A(\valid_counter[27] ),
    .B(_1683_),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _3699_ (.A(\valid_counter[26] ),
    .B(_1682_),
    .Y(_1690_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(_1683_),
    .B(_1690_),
    .Y(_0597_));
 sky130_fd_sc_hd__a31o_1 _3701_ (.A1(\valid_counter[24] ),
    .A2(\valid_counter[23] ),
    .A3(_1680_),
    .B1(\valid_counter[25] ),
    .X(_1691_));
 sky130_fd_sc_hd__and2b_1 _3702_ (.A_N(_1682_),
    .B(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__clkbuf_1 _3703_ (.A(_1692_),
    .X(_0596_));
 sky130_fd_sc_hd__xor2_1 _3704_ (.A(\valid_counter[24] ),
    .B(_1681_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _3705_ (.A(\valid_counter[23] ),
    .B(_1680_),
    .Y(_1693_));
 sky130_fd_sc_hd__nor2_1 _3706_ (.A(_1681_),
    .B(_1693_),
    .Y(_0594_));
 sky130_fd_sc_hd__a31o_1 _3707_ (.A1(\valid_counter[21] ),
    .A2(\valid_counter[20] ),
    .A3(_1678_),
    .B1(\valid_counter[22] ),
    .X(_1694_));
 sky130_fd_sc_hd__and2b_1 _3708_ (.A_N(_1680_),
    .B(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3709_ (.A(_1695_),
    .X(_0593_));
 sky130_fd_sc_hd__xor2_1 _3710_ (.A(\valid_counter[21] ),
    .B(_1679_),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _3711_ (.A(\valid_counter[20] ),
    .B(_1678_),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_1 _3712_ (.A(_1679_),
    .B(_1696_),
    .Y(_0591_));
 sky130_fd_sc_hd__a31o_1 _3713_ (.A1(\valid_counter[18] ),
    .A2(\valid_counter[17] ),
    .A3(_1676_),
    .B1(\valid_counter[19] ),
    .X(_1697_));
 sky130_fd_sc_hd__and2b_1 _3714_ (.A_N(_1678_),
    .B(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _3715_ (.A(_1698_),
    .X(_0590_));
 sky130_fd_sc_hd__xor2_1 _3716_ (.A(\valid_counter[18] ),
    .B(_1677_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _3717_ (.A(\valid_counter[17] ),
    .B(_1676_),
    .Y(_1699_));
 sky130_fd_sc_hd__nor2_1 _3718_ (.A(_1677_),
    .B(_1699_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(\valid_counter[15] ),
    .B(_1675_),
    .Y(_1700_));
 sky130_fd_sc_hd__xnor2_1 _3720_ (.A(\valid_counter[16] ),
    .B(_1700_),
    .Y(_0587_));
 sky130_fd_sc_hd__xor2_1 _3721_ (.A(\valid_counter[15] ),
    .B(_1675_),
    .X(_0586_));
 sky130_fd_sc_hd__xor2_1 _3722_ (.A(\valid_counter[14] ),
    .B(_1674_),
    .X(_0585_));
 sky130_fd_sc_hd__a31o_1 _3723_ (.A1(\valid_counter[12] ),
    .A2(\valid_counter[11] ),
    .A3(_1672_),
    .B1(\valid_counter[13] ),
    .X(_1701_));
 sky130_fd_sc_hd__and2b_1 _3724_ (.A_N(_1674_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _3725_ (.A(_1702_),
    .X(_0584_));
 sky130_fd_sc_hd__xor2_1 _3726_ (.A(\valid_counter[12] ),
    .B(_1673_),
    .X(_0583_));
 sky130_fd_sc_hd__nor2_1 _3727_ (.A(\valid_counter[11] ),
    .B(_1672_),
    .Y(_1703_));
 sky130_fd_sc_hd__nor2_1 _3728_ (.A(_1673_),
    .B(_1703_),
    .Y(_0582_));
 sky130_fd_sc_hd__a21oi_1 _3729_ (.A1(\valid_counter[9] ),
    .A2(_1671_),
    .B1(\valid_counter[10] ),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _3730_ (.A(_1672_),
    .B(_1704_),
    .Y(_0581_));
 sky130_fd_sc_hd__xor2_1 _3731_ (.A(\valid_counter[9] ),
    .B(_1671_),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _3732_ (.A(\valid_counter[8] ),
    .B(_1670_),
    .Y(_1705_));
 sky130_fd_sc_hd__nor2_1 _3733_ (.A(_1671_),
    .B(_1705_),
    .Y(_0579_));
 sky130_fd_sc_hd__a21oi_1 _3734_ (.A1(\valid_counter[6] ),
    .A2(_1669_),
    .B1(\valid_counter[7] ),
    .Y(_1706_));
 sky130_fd_sc_hd__nor2_1 _3735_ (.A(_1670_),
    .B(_1706_),
    .Y(_0578_));
 sky130_fd_sc_hd__xor2_1 _3736_ (.A(\valid_counter[6] ),
    .B(_1669_),
    .X(_0577_));
 sky130_fd_sc_hd__a31o_1 _3737_ (.A1(\valid_counter[4] ),
    .A2(\valid_counter[3] ),
    .A3(_1668_),
    .B1(\valid_counter[5] ),
    .X(_1707_));
 sky130_fd_sc_hd__and2b_1 _3738_ (.A_N(_1669_),
    .B(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _3739_ (.A(_1708_),
    .X(_0576_));
 sky130_fd_sc_hd__nand2_1 _3740_ (.A(\valid_counter[3] ),
    .B(_1668_),
    .Y(_1709_));
 sky130_fd_sc_hd__xnor2_1 _3741_ (.A(\valid_counter[4] ),
    .B(_1709_),
    .Y(_0575_));
 sky130_fd_sc_hd__or2_1 _3742_ (.A(\valid_counter[3] ),
    .B(_1668_),
    .X(_1710_));
 sky130_fd_sc_hd__and2_1 _3743_ (.A(_1709_),
    .B(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3744_ (.A(_1711_),
    .X(_0574_));
 sky130_fd_sc_hd__and3_1 _3745_ (.A(net10),
    .B(\valid_counter[1] ),
    .C(\valid_counter[0] ),
    .X(_1712_));
 sky130_fd_sc_hd__nor2_1 _3746_ (.A(\valid_counter[2] ),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2_1 _3747_ (.A(_1668_),
    .B(_1713_),
    .Y(_0573_));
 sky130_fd_sc_hd__a21oi_1 _3748_ (.A1(net10),
    .A2(\valid_counter[0] ),
    .B1(\valid_counter[1] ),
    .Y(_1714_));
 sky130_fd_sc_hd__nor2_1 _3749_ (.A(_1712_),
    .B(_1714_),
    .Y(_0572_));
 sky130_fd_sc_hd__xor2_1 _3750_ (.A(net10),
    .B(\valid_counter[0] ),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_2 _3751_ (.A(\col_operation[1] ),
    .X(_1715_));
 sky130_fd_sc_hd__clkbuf_2 _3752_ (.A(\col_operation[0] ),
    .X(_1716_));
 sky130_fd_sc_hd__and2_1 _3753_ (.A(_1715_),
    .B(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__and2_2 _3754_ (.A(\col_operation[3] ),
    .B(\col_operation[2] ),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__nand2_1 _3756_ (.A(_1717_),
    .B(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__a21o_1 _3757_ (.A1(_1079_),
    .A2(_1720_),
    .B1(_1427_),
    .X(_1721_));
 sky130_fd_sc_hd__and2_1 _3758_ (.A(_1079_),
    .B(_1099_),
    .X(_1722_));
 sky130_fd_sc_hd__and3b_2 _3759_ (.A_N(\col_operation[4] ),
    .B(_1715_),
    .C(_1716_),
    .X(_1723_));
 sky130_fd_sc_hd__and2_1 _3760_ (.A(_1718_),
    .B(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__buf_4 _3761_ (.A(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__buf_4 _3762_ (.A(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__buf_4 _3763_ (.A(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__buf_4 _3764_ (.A(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__a22o_1 _3765_ (.A1(\col_operation[4] ),
    .A2(_1721_),
    .B1(_1722_),
    .B2(_1728_),
    .X(_0570_));
 sky130_fd_sc_hd__nand2_1 _3766_ (.A(\col_operation[2] ),
    .B(_1717_),
    .Y(_1729_));
 sky130_fd_sc_hd__nor2_1 _3767_ (.A(_1427_),
    .B(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__o21a_1 _3768_ (.A1(\col_operation[3] ),
    .A2(_1730_),
    .B1(_1721_),
    .X(_0569_));
 sky130_fd_sc_hd__or2_1 _3769_ (.A(\col_operation[2] ),
    .B(_1717_),
    .X(_1731_));
 sky130_fd_sc_hd__a32o_1 _3770_ (.A1(_1729_),
    .A2(_1722_),
    .A3(_1731_),
    .B1(_1427_),
    .B2(\col_operation[2] ),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_2 _3771_ (.A(_1715_),
    .B(_1716_),
    .Y(_1732_));
 sky130_fd_sc_hd__o21ai_1 _3772_ (.A1(_1717_),
    .A2(_1732_),
    .B1(_1722_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21a_1 _3773_ (.A1(_1715_),
    .A2(_1099_),
    .B1(_1733_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _3774_ (.A0(_1722_),
    .A1(_1427_),
    .S(_1716_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _3775_ (.A(_1734_),
    .X(_0566_));
 sky130_fd_sc_hd__and3_1 _3776_ (.A(\col_input[5] ),
    .B(\col_input[4] ),
    .C(_1451_),
    .X(_1735_));
 sky130_fd_sc_hd__and4_1 _3777_ (.A(\col_input[8] ),
    .B(\col_input[7] ),
    .C(\col_input[6] ),
    .D(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__and4_1 _3778_ (.A(\col_input[11] ),
    .B(\col_input[10] ),
    .C(\col_input[9] ),
    .D(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__and4_1 _3779_ (.A(\col_input[14] ),
    .B(\col_input[13] ),
    .C(\col_input[12] ),
    .D(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__and3_1 _3780_ (.A(\col_input[16] ),
    .B(\col_input[15] ),
    .C(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__and2_1 _3781_ (.A(\col_input[17] ),
    .B(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__and3_1 _3782_ (.A(\col_input[19] ),
    .B(\col_input[18] ),
    .C(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__and2_1 _3783_ (.A(\col_input[20] ),
    .B(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__and3_1 _3784_ (.A(\col_input[22] ),
    .B(\col_input[21] ),
    .C(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__and2_1 _3785_ (.A(\col_input[23] ),
    .B(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__and3_1 _3786_ (.A(\col_input[25] ),
    .B(\col_input[24] ),
    .C(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__and2_1 _3787_ (.A(\col_input[26] ),
    .B(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__and3_1 _3788_ (.A(\col_input[28] ),
    .B(\col_input[27] ),
    .C(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__and2_1 _3789_ (.A(\col_input[29] ),
    .B(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a21oi_1 _3790_ (.A1(\col_input[30] ),
    .A2(_1748_),
    .B1(_1097_),
    .Y(_0565_));
 sky130_fd_sc_hd__xor2_1 _3791_ (.A(\col_input[30] ),
    .B(_1748_),
    .X(_0564_));
 sky130_fd_sc_hd__xor2_1 _3792_ (.A(\col_input[29] ),
    .B(_1747_),
    .X(_0563_));
 sky130_fd_sc_hd__a21oi_1 _3793_ (.A1(\col_input[27] ),
    .A2(_1746_),
    .B1(\col_input[28] ),
    .Y(_1749_));
 sky130_fd_sc_hd__nor2_1 _3794_ (.A(_1747_),
    .B(_1749_),
    .Y(_0562_));
 sky130_fd_sc_hd__xor2_1 _3795_ (.A(\col_input[27] ),
    .B(_1746_),
    .X(_0561_));
 sky130_fd_sc_hd__nor2_1 _3796_ (.A(\col_input[26] ),
    .B(_1745_),
    .Y(_1750_));
 sky130_fd_sc_hd__nor2_1 _3797_ (.A(_1746_),
    .B(_1750_),
    .Y(_0560_));
 sky130_fd_sc_hd__a21oi_1 _3798_ (.A1(\col_input[24] ),
    .A2(_1744_),
    .B1(\col_input[25] ),
    .Y(_1751_));
 sky130_fd_sc_hd__nor2_1 _3799_ (.A(_1745_),
    .B(_1751_),
    .Y(_0559_));
 sky130_fd_sc_hd__xor2_1 _3800_ (.A(\col_input[24] ),
    .B(_1744_),
    .X(_0558_));
 sky130_fd_sc_hd__xor2_1 _3801_ (.A(\col_input[23] ),
    .B(_1743_),
    .X(_0557_));
 sky130_fd_sc_hd__a31o_1 _3802_ (.A1(\col_input[21] ),
    .A2(\col_input[20] ),
    .A3(_1741_),
    .B1(\col_input[22] ),
    .X(_1752_));
 sky130_fd_sc_hd__and2b_1 _3803_ (.A_N(_1743_),
    .B(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__clkbuf_1 _3804_ (.A(_1753_),
    .X(_0556_));
 sky130_fd_sc_hd__xor2_1 _3805_ (.A(\col_input[21] ),
    .B(_1742_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _3806_ (.A(\col_input[20] ),
    .B(_1741_),
    .Y(_1754_));
 sky130_fd_sc_hd__nor2_1 _3807_ (.A(_1742_),
    .B(_1754_),
    .Y(_0554_));
 sky130_fd_sc_hd__a21oi_1 _3808_ (.A1(\col_input[18] ),
    .A2(_1740_),
    .B1(\col_input[19] ),
    .Y(_1755_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(_1741_),
    .B(_1755_),
    .Y(_0553_));
 sky130_fd_sc_hd__xor2_1 _3810_ (.A(\col_input[18] ),
    .B(_1740_),
    .X(_0552_));
 sky130_fd_sc_hd__nor2_1 _3811_ (.A(\col_input[17] ),
    .B(_1739_),
    .Y(_1756_));
 sky130_fd_sc_hd__nor2_1 _3812_ (.A(_1740_),
    .B(_1756_),
    .Y(_0551_));
 sky130_fd_sc_hd__a21oi_1 _3813_ (.A1(\col_input[15] ),
    .A2(_1738_),
    .B1(\col_input[16] ),
    .Y(_1757_));
 sky130_fd_sc_hd__nor2_1 _3814_ (.A(_1739_),
    .B(_1757_),
    .Y(_0550_));
 sky130_fd_sc_hd__xor2_1 _3815_ (.A(\col_input[15] ),
    .B(_1738_),
    .X(_0549_));
 sky130_fd_sc_hd__and3_1 _3816_ (.A(\col_input[13] ),
    .B(\col_input[12] ),
    .C(_1737_),
    .X(_1758_));
 sky130_fd_sc_hd__xor2_1 _3817_ (.A(\col_input[14] ),
    .B(_1758_),
    .X(_0548_));
 sky130_fd_sc_hd__a21oi_1 _3818_ (.A1(\col_input[12] ),
    .A2(_1737_),
    .B1(\col_input[13] ),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2_1 _3819_ (.A(_1758_),
    .B(_1759_),
    .Y(_0547_));
 sky130_fd_sc_hd__xor2_1 _3820_ (.A(\col_input[12] ),
    .B(_1737_),
    .X(_0546_));
 sky130_fd_sc_hd__nand3_1 _3821_ (.A(\col_input[10] ),
    .B(\col_input[9] ),
    .C(_1736_),
    .Y(_1760_));
 sky130_fd_sc_hd__xnor2_1 _3822_ (.A(\col_input[11] ),
    .B(_1760_),
    .Y(_0545_));
 sky130_fd_sc_hd__a21o_1 _3823_ (.A1(\col_input[9] ),
    .A2(_1736_),
    .B1(\col_input[10] ),
    .X(_1761_));
 sky130_fd_sc_hd__and2_1 _3824_ (.A(_1760_),
    .B(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__clkbuf_1 _3825_ (.A(_1762_),
    .X(_0544_));
 sky130_fd_sc_hd__xor2_1 _3826_ (.A(\col_input[9] ),
    .B(_1736_),
    .X(_0543_));
 sky130_fd_sc_hd__a31o_1 _3827_ (.A1(\col_input[7] ),
    .A2(\col_input[6] ),
    .A3(_1735_),
    .B1(\col_input[8] ),
    .X(_1763_));
 sky130_fd_sc_hd__and2b_1 _3828_ (.A_N(_1736_),
    .B(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3829_ (.A(_1764_),
    .X(_0542_));
 sky130_fd_sc_hd__and2_1 _3830_ (.A(\col_input[6] ),
    .B(_1735_),
    .X(_1765_));
 sky130_fd_sc_hd__xor2_1 _3831_ (.A(\col_input[7] ),
    .B(_1765_),
    .X(_0541_));
 sky130_fd_sc_hd__nor2_1 _3832_ (.A(\col_input[6] ),
    .B(_1735_),
    .Y(_1766_));
 sky130_fd_sc_hd__nor2_1 _3833_ (.A(_1765_),
    .B(_1766_),
    .Y(_0540_));
 sky130_fd_sc_hd__and2_1 _3834_ (.A(\col_input[4] ),
    .B(_1451_),
    .X(_1767_));
 sky130_fd_sc_hd__nor2_1 _3835_ (.A(\col_input[5] ),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__nor2_1 _3836_ (.A(_1735_),
    .B(_1768_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_1 _3837_ (.A(_1071_),
    .B(_1076_),
    .Y(_1769_));
 sky130_fd_sc_hd__a2bb2o_1 _3838_ (.A1_N(\col_input[4] ),
    .A2_N(_1451_),
    .B1(_1439_),
    .B2(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__nor2_1 _3839_ (.A(_1767_),
    .B(_1770_),
    .Y(_0538_));
 sky130_fd_sc_hd__nor2_1 _3840_ (.A(_1494_),
    .B(_1449_),
    .Y(_1771_));
 sky130_fd_sc_hd__xor2_1 _3841_ (.A(_1077_),
    .B(_1771_),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_1 _3842_ (.A(_1494_),
    .B(_1449_),
    .Y(_1772_));
 sky130_fd_sc_hd__and2b_1 _3843_ (.A_N(_1771_),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _3844_ (.A(_1773_),
    .X(_0536_));
 sky130_fd_sc_hd__nand2_1 _3845_ (.A(\col_input[0] ),
    .B(_1099_),
    .Y(_1774_));
 sky130_fd_sc_hd__xnor2_1 _3846_ (.A(\col_input[1] ),
    .B(_1774_),
    .Y(_0535_));
 sky130_fd_sc_hd__xnor2_1 _3847_ (.A(\col_input[0] ),
    .B(_1427_),
    .Y(_0534_));
 sky130_fd_sc_hd__clkbuf_4 _3848_ (.A(_1723_),
    .X(_1775_));
 sky130_fd_sc_hd__nor2_1 _3849_ (.A(\col_operation[3] ),
    .B(\col_operation[2] ),
    .Y(_1776_));
 sky130_fd_sc_hd__clkbuf_4 _3850_ (.A(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__nor2_1 _3851_ (.A(\col_operation[4] ),
    .B(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__nor3b_1 _3852_ (.A(\col_operation[3] ),
    .B(\col_operation[2] ),
    .C_N(\col_operation[4] ),
    .Y(_1779_));
 sky130_fd_sc_hd__clkbuf_4 _3853_ (.A(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__or3_1 _3854_ (.A(_1775_),
    .B(_1778_),
    .C(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__buf_4 _3855_ (.A(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__nor3b_1 _3856_ (.A(\col_operation[4] ),
    .B(_1715_),
    .C_N(_1716_),
    .Y(_1783_));
 sky130_fd_sc_hd__and2_1 _3857_ (.A(_1718_),
    .B(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__buf_4 _3858_ (.A(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__buf_4 _3859_ (.A(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__and3b_2 _3860_ (.A_N(_1716_),
    .B(_1780_),
    .C(_1715_),
    .X(_1787_));
 sky130_fd_sc_hd__buf_4 _3861_ (.A(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__and2_1 _3862_ (.A(_1723_),
    .B(_1776_),
    .X(_1789_));
 sky130_fd_sc_hd__buf_4 _3863_ (.A(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__and2_4 _3864_ (.A(_1717_),
    .B(_1780_),
    .X(_1791_));
 sky130_fd_sc_hd__a22o_1 _3865_ (.A1(\second_row[1][0] ),
    .A2(_1790_),
    .B1(_1791_),
    .B2(\second_row[17][0] ),
    .X(_1792_));
 sky130_fd_sc_hd__nor3_4 _3866_ (.A(_1775_),
    .B(_1778_),
    .C(_1780_),
    .Y(_1793_));
 sky130_fd_sc_hd__a211o_1 _3867_ (.A1(\second_row[16][0] ),
    .A2(_1788_),
    .B1(_1792_),
    .C1(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__and2b_1 _3868_ (.A_N(\col_operation[2] ),
    .B(\col_operation[3] ),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_4 _3869_ (.A(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__and2_1 _3870_ (.A(_1723_),
    .B(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__buf_4 _3871_ (.A(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_4 _3872_ (.A(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__nor3b_1 _3873_ (.A(\col_operation[4] ),
    .B(_1716_),
    .C_N(\col_operation[1] ),
    .Y(_1800_));
 sky130_fd_sc_hd__buf_2 _3874_ (.A(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__and2_2 _3875_ (.A(_1801_),
    .B(_1796_),
    .X(_1802_));
 sky130_fd_sc_hd__buf_4 _3876_ (.A(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__buf_4 _3877_ (.A(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__a22o_1 _3878_ (.A1(\second_row[9][0] ),
    .A2(_1799_),
    .B1(_1804_),
    .B2(\second_row[8][0] ),
    .X(_1805_));
 sky130_fd_sc_hd__a211o_1 _3879_ (.A1(\second_row[11][0] ),
    .A2(_1786_),
    .B1(_1794_),
    .C1(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__and3b_1 _3880_ (.A_N(_1715_),
    .B(_1716_),
    .C(_1780_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_4 _3881_ (.A(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__and2_1 _3882_ (.A(_1732_),
    .B(_1779_),
    .X(_1809_));
 sky130_fd_sc_hd__buf_4 _3883_ (.A(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__a22o_1 _3884_ (.A1(\second_row[13][0] ),
    .A2(_1725_),
    .B1(_1810_),
    .B2(\second_row[14][0] ),
    .X(_1811_));
 sky130_fd_sc_hd__and2_1 _3885_ (.A(_1783_),
    .B(_1796_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_4 _3886_ (.A(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__nor3_1 _3887_ (.A(\col_operation[4] ),
    .B(_1715_),
    .C(\col_operation[0] ),
    .Y(_1814_));
 sky130_fd_sc_hd__clkbuf_4 _3888_ (.A(_1814_),
    .X(_1815_));
 sky130_fd_sc_hd__and2_1 _3889_ (.A(_1718_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__buf_4 _3890_ (.A(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__and2_1 _3891_ (.A(_1718_),
    .B(_1801_),
    .X(_1818_));
 sky130_fd_sc_hd__buf_4 _3892_ (.A(_1818_),
    .X(_1819_));
 sky130_fd_sc_hd__and2b_1 _3893_ (.A_N(\col_operation[3] ),
    .B(\col_operation[2] ),
    .X(_1820_));
 sky130_fd_sc_hd__and2_1 _3894_ (.A(_1820_),
    .B(_1783_),
    .X(_1821_));
 sky130_fd_sc_hd__buf_4 _3895_ (.A(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__a22o_1 _3896_ (.A1(\second_row[12][0] ),
    .A2(_1819_),
    .B1(_1822_),
    .B2(\second_row[3][0] ),
    .X(_1823_));
 sky130_fd_sc_hd__a221o_1 _3897_ (.A1(\second_row[7][0] ),
    .A2(_1813_),
    .B1(_1817_),
    .B2(\second_row[10][0] ),
    .C1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__and2_1 _3898_ (.A(_1723_),
    .B(_1820_),
    .X(_1825_));
 sky130_fd_sc_hd__buf_4 _3899_ (.A(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__and2_1 _3900_ (.A(_1795_),
    .B(_1814_),
    .X(_1827_));
 sky130_fd_sc_hd__buf_4 _3901_ (.A(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__buf_4 _3902_ (.A(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__and2_1 _3903_ (.A(_1820_),
    .B(_1800_),
    .X(_1830_));
 sky130_fd_sc_hd__buf_4 _3904_ (.A(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__and2_1 _3905_ (.A(_1820_),
    .B(_1815_),
    .X(_1832_));
 sky130_fd_sc_hd__clkbuf_4 _3906_ (.A(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__a22o_1 _3907_ (.A1(\second_row[4][0] ),
    .A2(_1831_),
    .B1(_1833_),
    .B2(\second_row[2][0] ),
    .X(_1834_));
 sky130_fd_sc_hd__a221o_1 _3908_ (.A1(\second_row[5][0] ),
    .A2(_1826_),
    .B1(_1829_),
    .B2(\second_row[6][0] ),
    .C1(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__a2111o_2 _3909_ (.A1(\second_row[15][0] ),
    .A2(_1808_),
    .B1(_1811_),
    .C1(_1824_),
    .D1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__a22o_1 _3910_ (.A1(\first_row[6][0] ),
    .A2(_1826_),
    .B1(_1819_),
    .B2(\first_row[13][0] ),
    .X(_1837_));
 sky130_fd_sc_hd__a221o_1 _3911_ (.A1(\first_row[10][0] ),
    .A2(_1798_),
    .B1(_1817_),
    .B2(\first_row[11][0] ),
    .C1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__and3b_1 _3912_ (.A_N(_1716_),
    .B(_1777_),
    .C(_1715_),
    .X(_1839_));
 sky130_fd_sc_hd__or3_2 _3913_ (.A(\col_operation[3] ),
    .B(\col_operation[2] ),
    .C(_1715_),
    .X(_1840_));
 sky130_fd_sc_hd__xor2_4 _3914_ (.A(\col_operation[4] ),
    .B(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__nor2_4 _3915_ (.A(_1839_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__a21o_1 _3916_ (.A1(\first_row[16][0] ),
    .A2(_1808_),
    .B1(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__a22o_1 _3917_ (.A1(\first_row[8][0] ),
    .A2(_1812_),
    .B1(_1822_),
    .B2(\first_row[4][0] ),
    .X(_1844_));
 sky130_fd_sc_hd__a22o_1 _3918_ (.A1(\first_row[17][0] ),
    .A2(_1787_),
    .B1(_1802_),
    .B2(\first_row[9][0] ),
    .X(_1845_));
 sky130_fd_sc_hd__and3_1 _3919_ (.A(\first_row[1][0] ),
    .B(_1777_),
    .C(_1801_),
    .X(_1846_));
 sky130_fd_sc_hd__and3_1 _3920_ (.A(\first_row[7][0] ),
    .B(_1796_),
    .C(_1815_),
    .X(_1847_));
 sky130_fd_sc_hd__and3_1 _3921_ (.A(\first_row[14][0] ),
    .B(_1719_),
    .C(_1775_),
    .X(_1848_));
 sky130_fd_sc_hd__a2111o_1 _3922_ (.A1(\first_row[2][0] ),
    .A2(_1789_),
    .B1(_1846_),
    .C1(_1847_),
    .D1(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__buf_2 _3923_ (.A(_1820_),
    .X(_1850_));
 sky130_fd_sc_hd__and3_1 _3924_ (.A(\first_row[5][0] ),
    .B(_1850_),
    .C(_1801_),
    .X(_1851_));
 sky130_fd_sc_hd__and3_1 _3925_ (.A(\first_row[15][0] ),
    .B(_1732_),
    .C(_1780_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_4 _3926_ (.A(_1783_),
    .X(_1853_));
 sky130_fd_sc_hd__and3_1 _3927_ (.A(\first_row[12][0] ),
    .B(_1719_),
    .C(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__a2111o_1 _3928_ (.A1(\first_row[3][0] ),
    .A2(_1833_),
    .B1(_1851_),
    .C1(_1852_),
    .D1(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__or4_2 _3929_ (.A(_1844_),
    .B(_1845_),
    .C(_1849_),
    .D(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__or2_4 _3930_ (.A(_1839_),
    .B(_1841_),
    .X(_1857_));
 sky130_fd_sc_hd__o32a_1 _3931_ (.A1(_1838_),
    .A2(_1843_),
    .A3(_1856_),
    .B1(_1857_),
    .B2(\first_row[0][0] ),
    .X(_1858_));
 sky130_fd_sc_hd__o221a_1 _3932_ (.A1(\second_row[0][0] ),
    .A2(_1782_),
    .B1(_1806_),
    .B2(_1836_),
    .C1(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__o22a_1 _3933_ (.A1(\second_row[0][0] ),
    .A2(_1782_),
    .B1(_1806_),
    .B2(_1836_),
    .X(_1860_));
 sky130_fd_sc_hd__nor2_1 _3934_ (.A(_1860_),
    .B(_1858_),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _3935_ (.A(_1859_),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__and2b_2 _3936_ (.A_N(\col_operation[4] ),
    .B(_1716_),
    .X(_1863_));
 sky130_fd_sc_hd__or2_1 _3937_ (.A(_1863_),
    .B(_1841_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_8 _3938_ (.A(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__nor2_8 _3939_ (.A(_1863_),
    .B(_1841_),
    .Y(_1866_));
 sky130_fd_sc_hd__and2_1 _3940_ (.A(_1776_),
    .B(_1800_),
    .X(_1867_));
 sky130_fd_sc_hd__buf_4 _3941_ (.A(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__a22o_1 _3942_ (.A1(\second_row[14][0] ),
    .A2(_1819_),
    .B1(_1868_),
    .B2(\second_row[2][0] ),
    .X(_1869_));
 sky130_fd_sc_hd__a22o_1 _3943_ (.A1(\second_row[11][0] ),
    .A2(_1798_),
    .B1(_1785_),
    .B2(\second_row[13][0] ),
    .X(_1870_));
 sky130_fd_sc_hd__a22o_1 _3944_ (.A1(\second_row[6][0] ),
    .A2(_1831_),
    .B1(_1803_),
    .B2(\second_row[10][0] ),
    .X(_1871_));
 sky130_fd_sc_hd__or4_4 _3945_ (.A(_1866_),
    .B(_1869_),
    .C(_1870_),
    .D(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__and3_1 _3946_ (.A(\second_row[7][0] ),
    .B(_1775_),
    .C(_1850_),
    .X(_1873_));
 sky130_fd_sc_hd__and3_1 _3947_ (.A(\second_row[16][0] ),
    .B(_1732_),
    .C(_1780_),
    .X(_1874_));
 sky130_fd_sc_hd__a221o_1 _3948_ (.A1(\second_row[15][0] ),
    .A2(_1725_),
    .B1(_1808_),
    .B2(\second_row[17][0] ),
    .C1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__a22o_1 _3949_ (.A1(\second_row[12][0] ),
    .A2(_1817_),
    .B1(_1833_),
    .B2(\second_row[4][0] ),
    .X(_1876_));
 sky130_fd_sc_hd__and2_4 _3950_ (.A(_1777_),
    .B(_1853_),
    .X(_1877_));
 sky130_fd_sc_hd__a22o_1 _3951_ (.A1(\second_row[3][0] ),
    .A2(_1790_),
    .B1(_1877_),
    .B2(\second_row[1][0] ),
    .X(_1878_));
 sky130_fd_sc_hd__a22o_1 _3952_ (.A1(\second_row[9][0] ),
    .A2(_1813_),
    .B1(_1822_),
    .B2(\second_row[5][0] ),
    .X(_1879_));
 sky130_fd_sc_hd__a211o_1 _3953_ (.A1(\second_row[8][0] ),
    .A2(_1828_),
    .B1(_1878_),
    .C1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__or4_2 _3954_ (.A(_1873_),
    .B(_1875_),
    .C(_1876_),
    .D(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__and3_1 _3955_ (.A(\third_row[15][0] ),
    .B(_1732_),
    .C(_1780_),
    .X(_1882_));
 sky130_fd_sc_hd__a221o_1 _3956_ (.A1(\third_row[14][0] ),
    .A2(_1725_),
    .B1(_1808_),
    .B2(\third_row[16][0] ),
    .C1(_1882_),
    .X(_1883_));
 sky130_fd_sc_hd__a221o_1 _3957_ (.A1(\third_row[2][0] ),
    .A2(_1790_),
    .B1(_1829_),
    .B2(\third_row[7][0] ),
    .C1(_1842_),
    .X(_1884_));
 sky130_fd_sc_hd__and3_1 _3958_ (.A(\third_row[3][0] ),
    .B(_1850_),
    .C(_1815_),
    .X(_1885_));
 sky130_fd_sc_hd__and3_1 _3959_ (.A(\third_row[1][0] ),
    .B(_1777_),
    .C(_1801_),
    .X(_1886_));
 sky130_fd_sc_hd__and3_1 _3960_ (.A(\third_row[11][0] ),
    .B(_1719_),
    .C(_1815_),
    .X(_1887_));
 sky130_fd_sc_hd__a2111o_1 _3961_ (.A1(\third_row[17][0] ),
    .A2(_1787_),
    .B1(_1885_),
    .C1(_1886_),
    .D1(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__and3_1 _3962_ (.A(\third_row[4][0] ),
    .B(_1850_),
    .C(_1853_),
    .X(_1889_));
 sky130_fd_sc_hd__a221o_1 _3963_ (.A1(\third_row[12][0] ),
    .A2(_1785_),
    .B1(_1803_),
    .B2(\third_row[9][0] ),
    .C1(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__and3_1 _3964_ (.A(\third_row[5][0] ),
    .B(_1850_),
    .C(_1801_),
    .X(_1891_));
 sky130_fd_sc_hd__and3_1 _3965_ (.A(\third_row[13][0] ),
    .B(_1719_),
    .C(_1801_),
    .X(_1892_));
 sky130_fd_sc_hd__and3_1 _3966_ (.A(\third_row[6][0] ),
    .B(_1775_),
    .C(_1850_),
    .X(_1893_));
 sky130_fd_sc_hd__a2111o_1 _3967_ (.A1(\third_row[8][0] ),
    .A2(_1813_),
    .B1(_1891_),
    .C1(_1892_),
    .D1(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__a2111o_1 _3968_ (.A1(\third_row[10][0] ),
    .A2(_1798_),
    .B1(_1888_),
    .C1(_1890_),
    .D1(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__o32a_2 _3969_ (.A1(_1883_),
    .A2(_1884_),
    .A3(_1895_),
    .B1(_1857_),
    .B2(\third_row[0][0] ),
    .X(_1896_));
 sky130_fd_sc_hd__o221a_1 _3970_ (.A1(\second_row[0][0] ),
    .A2(_1865_),
    .B1(_1872_),
    .B2(_1881_),
    .C1(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__o22a_1 _3971_ (.A1(\second_row[0][0] ),
    .A2(_1865_),
    .B1(_1872_),
    .B2(_1881_),
    .X(_1898_));
 sky130_fd_sc_hd__nor2_1 _3972_ (.A(_1896_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__nor2_1 _3973_ (.A(_1897_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__and2_1 _3974_ (.A(_1862_),
    .B(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(_1862_),
    .B(_1900_),
    .Y(_1902_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_1901_),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__buf_4 _3977_ (.A(_1857_),
    .X(_1904_));
 sky130_fd_sc_hd__buf_4 _3978_ (.A(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__buf_4 _3979_ (.A(_1826_),
    .X(_1906_));
 sky130_fd_sc_hd__buf_4 _3980_ (.A(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_4 _3981_ (.A(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__buf_4 _3982_ (.A(_1804_),
    .X(_1909_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__buf_4 _3984_ (.A(_1819_),
    .X(_1911_));
 sky130_fd_sc_hd__buf_4 _3985_ (.A(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__buf_4 _3986_ (.A(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__buf_4 _3987_ (.A(_1822_),
    .X(_1914_));
 sky130_fd_sc_hd__clkbuf_4 _3988_ (.A(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__buf_4 _3989_ (.A(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__a22o_1 _3990_ (.A1(\second_row[13][6] ),
    .A2(_1913_),
    .B1(_1916_),
    .B2(\second_row[4][6] ),
    .X(_1917_));
 sky130_fd_sc_hd__a221o_1 _3991_ (.A1(\second_row[6][6] ),
    .A2(_1908_),
    .B1(_1910_),
    .B2(\second_row[9][6] ),
    .C1(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__buf_4 _3992_ (.A(_1842_),
    .X(_1919_));
 sky130_fd_sc_hd__buf_4 _3993_ (.A(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__buf_4 _3994_ (.A(_1829_),
    .X(_1921_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__buf_4 _3996_ (.A(_1810_),
    .X(_1923_));
 sky130_fd_sc_hd__buf_4 _3997_ (.A(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__clkbuf_4 _3998_ (.A(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__buf_4 _3999_ (.A(_1817_),
    .X(_1926_));
 sky130_fd_sc_hd__buf_4 _4000_ (.A(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__clkbuf_4 _4001_ (.A(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__buf_4 _4002_ (.A(_1868_),
    .X(_1929_));
 sky130_fd_sc_hd__buf_4 _4003_ (.A(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__a22o_1 _4004_ (.A1(\second_row[11][6] ),
    .A2(_1928_),
    .B1(_1930_),
    .B2(\second_row[1][6] ),
    .X(_1931_));
 sky130_fd_sc_hd__a221o_1 _4005_ (.A1(\second_row[7][6] ),
    .A2(_1922_),
    .B1(_1925_),
    .B2(\second_row[15][6] ),
    .C1(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__buf_4 _4006_ (.A(_1808_),
    .X(_1933_));
 sky130_fd_sc_hd__buf_4 _4007_ (.A(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_4 _4008_ (.A(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__clkbuf_4 _4009_ (.A(_1790_),
    .X(_1936_));
 sky130_fd_sc_hd__buf_4 _4010_ (.A(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__clkbuf_4 _4011_ (.A(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__buf_4 _4012_ (.A(_1833_),
    .X(_1939_));
 sky130_fd_sc_hd__buf_4 _4013_ (.A(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_4 _4014_ (.A(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__a22o_1 _4015_ (.A1(\second_row[2][6] ),
    .A2(_1938_),
    .B1(_1941_),
    .B2(\second_row[3][6] ),
    .X(_1942_));
 sky130_fd_sc_hd__buf_4 _4016_ (.A(_1788_),
    .X(_1943_));
 sky130_fd_sc_hd__buf_4 _4017_ (.A(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__buf_4 _4018_ (.A(_1799_),
    .X(_1945_));
 sky130_fd_sc_hd__buf_4 _4019_ (.A(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__a22o_1 _4020_ (.A1(\second_row[17][6] ),
    .A2(_1944_),
    .B1(_1946_),
    .B2(\second_row[10][6] ),
    .X(_1947_));
 sky130_fd_sc_hd__a211o_1 _4021_ (.A1(\second_row[16][6] ),
    .A2(_1935_),
    .B1(_1942_),
    .C1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__buf_4 _4022_ (.A(_1786_),
    .X(_1949_));
 sky130_fd_sc_hd__buf_4 _4023_ (.A(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__buf_4 _4024_ (.A(_1831_),
    .X(_1951_));
 sky130_fd_sc_hd__clkbuf_4 _4025_ (.A(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__buf_4 _4026_ (.A(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__buf_4 _4027_ (.A(_1813_),
    .X(_1954_));
 sky130_fd_sc_hd__buf_4 _4028_ (.A(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__buf_4 _4029_ (.A(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__a22o_1 _4030_ (.A1(\second_row[5][6] ),
    .A2(_1953_),
    .B1(_1956_),
    .B2(\second_row[8][6] ),
    .X(_1957_));
 sky130_fd_sc_hd__a221o_1 _4031_ (.A1(\second_row[14][6] ),
    .A2(_1728_),
    .B1(_1950_),
    .B2(\second_row[12][6] ),
    .C1(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__or4_1 _4032_ (.A(_1920_),
    .B(_1932_),
    .C(_1948_),
    .D(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__o22a_1 _4033_ (.A1(\second_row[0][6] ),
    .A2(_1905_),
    .B1(_1918_),
    .B2(_1959_),
    .X(_1960_));
 sky130_fd_sc_hd__a22o_1 _4034_ (.A1(\second_row[15][3] ),
    .A2(_1925_),
    .B1(_1941_),
    .B2(\second_row[3][3] ),
    .X(_1961_));
 sky130_fd_sc_hd__a221o_1 _4035_ (.A1(\second_row[14][3] ),
    .A2(_1728_),
    .B1(_1946_),
    .B2(\second_row[10][3] ),
    .C1(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__a211o_1 _4036_ (.A1(\second_row[16][3] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__a22o_1 _4037_ (.A1(\second_row[13][3] ),
    .A2(_1913_),
    .B1(_1928_),
    .B2(\second_row[11][3] ),
    .X(_1964_));
 sky130_fd_sc_hd__a221o_1 _4038_ (.A1(\second_row[6][3] ),
    .A2(_1908_),
    .B1(_1922_),
    .B2(\second_row[7][3] ),
    .C1(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__a22o_1 _4039_ (.A1(\second_row[2][3] ),
    .A2(_1938_),
    .B1(_1930_),
    .B2(\second_row[1][3] ),
    .X(_1966_));
 sky130_fd_sc_hd__a221o_1 _4040_ (.A1(\second_row[8][3] ),
    .A2(_1956_),
    .B1(_1950_),
    .B2(\second_row[12][3] ),
    .C1(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__a22o_1 _4041_ (.A1(\second_row[5][3] ),
    .A2(_1953_),
    .B1(_1916_),
    .B2(\second_row[4][3] ),
    .X(_1968_));
 sky130_fd_sc_hd__a221o_1 _4042_ (.A1(\second_row[17][3] ),
    .A2(_1944_),
    .B1(_1910_),
    .B2(\second_row[9][3] ),
    .C1(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__or3_2 _4043_ (.A(_1965_),
    .B(_1967_),
    .C(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__o22a_1 _4044_ (.A1(\second_row[0][3] ),
    .A2(_1905_),
    .B1(_1963_),
    .B2(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__a22o_1 _4045_ (.A1(\second_row[14][2] ),
    .A2(_1727_),
    .B1(_1930_),
    .B2(\second_row[1][2] ),
    .X(_1972_));
 sky130_fd_sc_hd__a221o_1 _4046_ (.A1(\second_row[5][2] ),
    .A2(_1953_),
    .B1(_1910_),
    .B2(\second_row[9][2] ),
    .C1(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__a211o_1 _4047_ (.A1(\second_row[16][2] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_1973_),
    .X(_1974_));
 sky130_fd_sc_hd__a22o_1 _4048_ (.A1(\second_row[11][2] ),
    .A2(_1928_),
    .B1(_1922_),
    .B2(\second_row[7][2] ),
    .X(_1975_));
 sky130_fd_sc_hd__a221o_1 _4049_ (.A1(\second_row[10][2] ),
    .A2(_1946_),
    .B1(_1950_),
    .B2(\second_row[12][2] ),
    .C1(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a22o_1 _4050_ (.A1(\second_row[2][2] ),
    .A2(_1938_),
    .B1(_1912_),
    .B2(\second_row[13][2] ),
    .X(_1977_));
 sky130_fd_sc_hd__a221o_1 _4051_ (.A1(\second_row[17][2] ),
    .A2(_1944_),
    .B1(_1956_),
    .B2(\second_row[8][2] ),
    .C1(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__a22o_1 _4052_ (.A1(\second_row[6][2] ),
    .A2(_1908_),
    .B1(_1941_),
    .B2(\second_row[3][2] ),
    .X(_1979_));
 sky130_fd_sc_hd__a221o_1 _4053_ (.A1(\second_row[4][2] ),
    .A2(_1916_),
    .B1(_1925_),
    .B2(\second_row[15][2] ),
    .C1(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__or3_1 _4054_ (.A(_1976_),
    .B(_1978_),
    .C(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__o22a_1 _4055_ (.A1(\second_row[0][2] ),
    .A2(_1905_),
    .B1(_1974_),
    .B2(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__nor2_1 _4056_ (.A(\second_row[0][1] ),
    .B(_1905_),
    .Y(_1983_));
 sky130_fd_sc_hd__a22o_1 _4057_ (.A1(\second_row[8][1] ),
    .A2(_1956_),
    .B1(_1910_),
    .B2(\second_row[9][1] ),
    .X(_1984_));
 sky130_fd_sc_hd__a221o_1 _4058_ (.A1(\second_row[14][1] ),
    .A2(_1728_),
    .B1(_1913_),
    .B2(\second_row[13][1] ),
    .C1(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__a22o_1 _4059_ (.A1(\second_row[6][1] ),
    .A2(_1907_),
    .B1(_1949_),
    .B2(\second_row[12][1] ),
    .X(_1986_));
 sky130_fd_sc_hd__a221o_1 _4060_ (.A1(\second_row[5][1] ),
    .A2(_1952_),
    .B1(_1916_),
    .B2(\second_row[4][1] ),
    .C1(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__a22o_1 _4061_ (.A1(\second_row[2][1] ),
    .A2(_1937_),
    .B1(_1927_),
    .B2(\second_row[11][1] ),
    .X(_1988_));
 sky130_fd_sc_hd__a22o_1 _4062_ (.A1(\second_row[7][1] ),
    .A2(_1921_),
    .B1(_1924_),
    .B2(\second_row[15][1] ),
    .X(_1989_));
 sky130_fd_sc_hd__a211o_1 _4063_ (.A1(\second_row[16][1] ),
    .A2(_1934_),
    .B1(_1988_),
    .C1(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__a22o_1 _4064_ (.A1(\second_row[10][1] ),
    .A2(_1945_),
    .B1(_1930_),
    .B2(\second_row[1][1] ),
    .X(_1991_));
 sky130_fd_sc_hd__a221o_1 _4065_ (.A1(\second_row[17][1] ),
    .A2(_1944_),
    .B1(_1941_),
    .B2(\second_row[3][1] ),
    .C1(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__or4_1 _4066_ (.A(_1920_),
    .B(_1987_),
    .C(_1990_),
    .D(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__nor2_1 _4067_ (.A(_1985_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(\second_row[8][0] ),
    .A2(_1955_),
    .B1(_1909_),
    .B2(\second_row[9][0] ),
    .X(_1995_));
 sky130_fd_sc_hd__a22o_1 _4069_ (.A1(\second_row[13][0] ),
    .A2(_1912_),
    .B1(_1945_),
    .B2(\second_row[10][0] ),
    .X(_1996_));
 sky130_fd_sc_hd__a221o_1 _4070_ (.A1(\second_row[6][0] ),
    .A2(_1907_),
    .B1(_1952_),
    .B2(\second_row[5][0] ),
    .C1(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__a22o_1 _4071_ (.A1(\second_row[14][0] ),
    .A2(_1727_),
    .B1(_1915_),
    .B2(\second_row[4][0] ),
    .X(_1998_));
 sky130_fd_sc_hd__a22o_1 _4072_ (.A1(\second_row[17][0] ),
    .A2(_1943_),
    .B1(_1940_),
    .B2(\second_row[3][0] ),
    .X(_1999_));
 sky130_fd_sc_hd__a221o_1 _4073_ (.A1(\second_row[2][0] ),
    .A2(_1937_),
    .B1(_1921_),
    .B2(\second_row[7][0] ),
    .C1(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__a221o_1 _4074_ (.A1(\second_row[11][0] ),
    .A2(_1926_),
    .B1(_1929_),
    .B2(\second_row[1][0] ),
    .C1(_1919_),
    .X(_2001_));
 sky130_fd_sc_hd__a221o_1 _4075_ (.A1(\second_row[16][0] ),
    .A2(_1933_),
    .B1(_1924_),
    .B2(\second_row[15][0] ),
    .C1(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__or4_1 _4076_ (.A(_1997_),
    .B(_1998_),
    .C(_2000_),
    .D(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__a211o_1 _4077_ (.A1(\second_row[12][0] ),
    .A2(_1950_),
    .B1(_1995_),
    .C1(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__o21ai_2 _4078_ (.A1(\second_row[0][0] ),
    .A2(_1905_),
    .B1(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__o21a_1 _4079_ (.A1(_1983_),
    .A2(_1994_),
    .B1(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__and2b_1 _4080_ (.A_N(_1982_),
    .B(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__and2b_2 _4081_ (.A_N(_1971_),
    .B(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__a22o_1 _4082_ (.A1(\second_row[5][4] ),
    .A2(_1953_),
    .B1(_1916_),
    .B2(\second_row[4][4] ),
    .X(_2009_));
 sky130_fd_sc_hd__a221o_2 _4083_ (.A1(\second_row[13][4] ),
    .A2(_1913_),
    .B1(_1950_),
    .B2(\second_row[12][4] ),
    .C1(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__a22o_1 _4084_ (.A1(\second_row[17][4] ),
    .A2(_1944_),
    .B1(_1922_),
    .B2(\second_row[7][4] ),
    .X(_2011_));
 sky130_fd_sc_hd__a221o_1 _4085_ (.A1(\second_row[2][4] ),
    .A2(_1938_),
    .B1(_1925_),
    .B2(\second_row[15][4] ),
    .C1(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__a22o_1 _4086_ (.A1(\second_row[10][4] ),
    .A2(_1946_),
    .B1(_1928_),
    .B2(\second_row[11][4] ),
    .X(_2013_));
 sky130_fd_sc_hd__a221o_1 _4087_ (.A1(\second_row[3][4] ),
    .A2(_1941_),
    .B1(_1930_),
    .B2(\second_row[1][4] ),
    .C1(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__a211o_1 _4088_ (.A1(\second_row[16][4] ),
    .A2(_1935_),
    .B1(_2012_),
    .C1(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__a22o_1 _4089_ (.A1(\second_row[8][4] ),
    .A2(_1956_),
    .B1(_1910_),
    .B2(\second_row[9][4] ),
    .X(_2016_));
 sky130_fd_sc_hd__a221o_1 _4090_ (.A1(\second_row[14][4] ),
    .A2(_1728_),
    .B1(_1908_),
    .B2(\second_row[6][4] ),
    .C1(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__or3_2 _4091_ (.A(_1920_),
    .B(_2015_),
    .C(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__o22ai_4 _4092_ (.A1(\second_row[0][4] ),
    .A2(_1905_),
    .B1(_2010_),
    .B2(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__a22o_1 _4093_ (.A1(\second_row[13][5] ),
    .A2(_1913_),
    .B1(_1950_),
    .B2(\second_row[12][5] ),
    .X(_2020_));
 sky130_fd_sc_hd__a221o_1 _4094_ (.A1(\second_row[5][5] ),
    .A2(_1953_),
    .B1(_1916_),
    .B2(\second_row[4][5] ),
    .C1(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__a22o_1 _4095_ (.A1(\second_row[17][5] ),
    .A2(_1944_),
    .B1(_1941_),
    .B2(\second_row[3][5] ),
    .X(_2022_));
 sky130_fd_sc_hd__a221o_1 _4096_ (.A1(\second_row[2][5] ),
    .A2(_1938_),
    .B1(_1928_),
    .B2(\second_row[11][5] ),
    .C1(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a22o_1 _4097_ (.A1(\second_row[7][5] ),
    .A2(_1922_),
    .B1(_1930_),
    .B2(\second_row[1][5] ),
    .X(_2024_));
 sky130_fd_sc_hd__a221o_1 _4098_ (.A1(\second_row[10][5] ),
    .A2(_1946_),
    .B1(_1925_),
    .B2(\second_row[15][5] ),
    .C1(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__a2111o_1 _4099_ (.A1(\second_row[16][5] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_2023_),
    .D1(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__a22o_1 _4100_ (.A1(\second_row[14][5] ),
    .A2(_1728_),
    .B1(_1908_),
    .B2(\second_row[6][5] ),
    .X(_2027_));
 sky130_fd_sc_hd__a221o_1 _4101_ (.A1(\second_row[8][5] ),
    .A2(_1956_),
    .B1(_1910_),
    .B2(\second_row[9][5] ),
    .C1(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__or3_1 _4102_ (.A(_2021_),
    .B(_2026_),
    .C(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__o21ai_1 _4103_ (.A1(\second_row[0][5] ),
    .A2(_1905_),
    .B1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__and3_1 _4104_ (.A(_2008_),
    .B(_2019_),
    .C(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__and2b_1 _4105_ (.A_N(_1960_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__a22o_1 _4106_ (.A1(\second_row[14][7] ),
    .A2(_1728_),
    .B1(_1938_),
    .B2(\second_row[2][7] ),
    .X(_2033_));
 sky130_fd_sc_hd__a221o_1 _4107_ (.A1(\second_row[8][7] ),
    .A2(_1956_),
    .B1(_1930_),
    .B2(\second_row[1][7] ),
    .C1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__a211o_1 _4108_ (.A1(\second_row[16][7] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__a22o_1 _4109_ (.A1(\second_row[17][7] ),
    .A2(_1944_),
    .B1(_1941_),
    .B2(\second_row[3][7] ),
    .X(_2036_));
 sky130_fd_sc_hd__a221o_1 _4110_ (.A1(\second_row[12][7] ),
    .A2(_1950_),
    .B1(_1925_),
    .B2(\second_row[15][7] ),
    .C1(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__a22o_1 _4111_ (.A1(\second_row[11][7] ),
    .A2(_1928_),
    .B1(_1922_),
    .B2(\second_row[7][7] ),
    .X(_2038_));
 sky130_fd_sc_hd__a221o_1 _4112_ (.A1(\second_row[5][7] ),
    .A2(_1953_),
    .B1(_1910_),
    .B2(\second_row[9][7] ),
    .C1(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(\second_row[13][7] ),
    .A2(_1913_),
    .B1(_1946_),
    .B2(\second_row[10][7] ),
    .X(_2040_));
 sky130_fd_sc_hd__a221o_1 _4114_ (.A1(\second_row[6][7] ),
    .A2(_1908_),
    .B1(_1916_),
    .B2(\second_row[4][7] ),
    .C1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__or3_1 _4115_ (.A(_2037_),
    .B(_2039_),
    .C(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__o22a_1 _4116_ (.A1(\second_row[0][7] ),
    .A2(_1905_),
    .B1(_2035_),
    .B2(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__xnor2_1 _4117_ (.A(_2032_),
    .B(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__nor2_1 _4118_ (.A(\first_row[0][7] ),
    .B(_1905_),
    .Y(_2045_));
 sky130_fd_sc_hd__a22o_1 _4119_ (.A1(\first_row[8][7] ),
    .A2(_1956_),
    .B1(_1946_),
    .B2(\first_row[10][7] ),
    .X(_2046_));
 sky130_fd_sc_hd__a221o_1 _4120_ (.A1(\first_row[6][7] ),
    .A2(_1908_),
    .B1(_1910_),
    .B2(\first_row[9][7] ),
    .C1(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__a22o_1 _4121_ (.A1(\first_row[5][7] ),
    .A2(_1953_),
    .B1(_1916_),
    .B2(\first_row[4][7] ),
    .X(_2048_));
 sky130_fd_sc_hd__a221o_1 _4122_ (.A1(\first_row[14][7] ),
    .A2(_1728_),
    .B1(_1950_),
    .B2(\first_row[12][7] ),
    .C1(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__a22o_1 _4123_ (.A1(\first_row[17][7] ),
    .A2(_1944_),
    .B1(_1930_),
    .B2(\first_row[1][7] ),
    .X(_2050_));
 sky130_fd_sc_hd__a221o_1 _4124_ (.A1(\first_row[13][7] ),
    .A2(_1913_),
    .B1(_1928_),
    .B2(\first_row[11][7] ),
    .C1(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__a22o_1 _4125_ (.A1(\first_row[2][7] ),
    .A2(_1938_),
    .B1(_1922_),
    .B2(\first_row[7][7] ),
    .X(_2052_));
 sky130_fd_sc_hd__a221o_1 _4126_ (.A1(\first_row[15][7] ),
    .A2(_1925_),
    .B1(_1941_),
    .B2(\first_row[3][7] ),
    .C1(_2052_),
    .X(_2053_));
 sky130_fd_sc_hd__a2111o_1 _4127_ (.A1(\first_row[16][7] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_2051_),
    .D1(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__nor3_1 _4128_ (.A(_2047_),
    .B(_2049_),
    .C(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__nor2_1 _4129_ (.A(\second_row[0][7] ),
    .B(_1782_),
    .Y(_2056_));
 sky130_fd_sc_hd__a22o_1 _4130_ (.A1(\second_row[7][7] ),
    .A2(_1955_),
    .B1(_1946_),
    .B2(\second_row[9][7] ),
    .X(_2057_));
 sky130_fd_sc_hd__a221o_1 _4131_ (.A1(\second_row[12][7] ),
    .A2(_1913_),
    .B1(_1910_),
    .B2(\second_row[8][7] ),
    .C1(_2057_),
    .X(_2058_));
 sky130_fd_sc_hd__a221o_1 _4132_ (.A1(\second_row[15][7] ),
    .A2(_1935_),
    .B1(_1922_),
    .B2(\second_row[6][7] ),
    .C1(_1793_),
    .X(_2059_));
 sky130_fd_sc_hd__or2_1 _4133_ (.A(_2058_),
    .B(_2059_),
    .X(_2060_));
 sky130_fd_sc_hd__a22o_1 _4134_ (.A1(\second_row[13][7] ),
    .A2(_1728_),
    .B1(_1938_),
    .B2(\second_row[1][7] ),
    .X(_2061_));
 sky130_fd_sc_hd__a22o_1 _4135_ (.A1(\second_row[3][7] ),
    .A2(_1915_),
    .B1(_1941_),
    .B2(\second_row[2][7] ),
    .X(_2062_));
 sky130_fd_sc_hd__a221o_1 _4136_ (.A1(\second_row[11][7] ),
    .A2(_1950_),
    .B1(_1925_),
    .B2(\second_row[14][7] ),
    .C1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__a22o_1 _4137_ (.A1(\second_row[5][7] ),
    .A2(_1908_),
    .B1(_1791_),
    .B2(\second_row[17][7] ),
    .X(_2064_));
 sky130_fd_sc_hd__a221o_1 _4138_ (.A1(\second_row[16][7] ),
    .A2(_1944_),
    .B1(_1928_),
    .B2(\second_row[10][7] ),
    .C1(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__a2111o_1 _4139_ (.A1(\second_row[4][7] ),
    .A2(_1953_),
    .B1(_2061_),
    .C1(_2063_),
    .D1(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__nor2_1 _4140_ (.A(_2060_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__o22a_1 _4141_ (.A1(_2045_),
    .A2(_2055_),
    .B1(_2056_),
    .B2(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__nor4_1 _4142_ (.A(_2045_),
    .B(_2055_),
    .C(_2056_),
    .D(_2067_),
    .Y(_2069_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(\first_row[0][5] ),
    .B(_1904_),
    .Y(_2070_));
 sky130_fd_sc_hd__a22o_1 _4144_ (.A1(\first_row[8][5] ),
    .A2(_1955_),
    .B1(_1945_),
    .B2(\first_row[10][5] ),
    .X(_2071_));
 sky130_fd_sc_hd__a221o_1 _4145_ (.A1(\first_row[6][5] ),
    .A2(_1907_),
    .B1(_1912_),
    .B2(\first_row[13][5] ),
    .C1(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__a22o_2 _4146_ (.A1(\first_row[5][5] ),
    .A2(_1952_),
    .B1(_1915_),
    .B2(\first_row[4][5] ),
    .X(_2073_));
 sky130_fd_sc_hd__a221o_1 _4147_ (.A1(\first_row[12][5] ),
    .A2(_1949_),
    .B1(_1909_),
    .B2(\first_row[9][5] ),
    .C1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__a22o_1 _4148_ (.A1(\first_row[11][5] ),
    .A2(_1926_),
    .B1(_1929_),
    .B2(\first_row[1][5] ),
    .X(_2075_));
 sky130_fd_sc_hd__a221o_1 _4149_ (.A1(\first_row[7][5] ),
    .A2(_1921_),
    .B1(_1924_),
    .B2(\first_row[15][5] ),
    .C1(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__a22o_1 _4150_ (.A1(\first_row[14][5] ),
    .A2(_1726_),
    .B1(_1943_),
    .B2(\first_row[17][5] ),
    .X(_2077_));
 sky130_fd_sc_hd__a221o_1 _4151_ (.A1(\first_row[2][5] ),
    .A2(_1937_),
    .B1(_1940_),
    .B2(\first_row[3][5] ),
    .C1(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__a2111o_1 _4152_ (.A1(\first_row[16][5] ),
    .A2(_1934_),
    .B1(_1919_),
    .C1(_2076_),
    .D1(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__nor3_1 _4153_ (.A(_2072_),
    .B(_2074_),
    .C(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__nor2_1 _4154_ (.A(\second_row[0][5] ),
    .B(_1782_),
    .Y(_2081_));
 sky130_fd_sc_hd__a22o_1 _4155_ (.A1(\second_row[12][5] ),
    .A2(_1912_),
    .B1(_1949_),
    .B2(\second_row[11][5] ),
    .X(_2082_));
 sky130_fd_sc_hd__a221o_1 _4156_ (.A1(\second_row[4][5] ),
    .A2(_1952_),
    .B1(_1925_),
    .B2(\second_row[14][5] ),
    .C1(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__a221o_1 _4157_ (.A1(\second_row[15][5] ),
    .A2(_1934_),
    .B1(_1909_),
    .B2(\second_row[8][5] ),
    .C1(_1793_),
    .X(_2084_));
 sky130_fd_sc_hd__a22o_1 _4158_ (.A1(\second_row[17][5] ),
    .A2(_1791_),
    .B1(_1940_),
    .B2(\second_row[2][5] ),
    .X(_2085_));
 sky130_fd_sc_hd__a22o_1 _4159_ (.A1(\second_row[16][5] ),
    .A2(_1943_),
    .B1(_1954_),
    .B2(\second_row[7][5] ),
    .X(_2086_));
 sky130_fd_sc_hd__a221o_1 _4160_ (.A1(\second_row[10][5] ),
    .A2(_1927_),
    .B1(_1921_),
    .B2(\second_row[6][5] ),
    .C1(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a22o_1 _4161_ (.A1(\second_row[9][5] ),
    .A2(_1945_),
    .B1(_1914_),
    .B2(\second_row[3][5] ),
    .X(_2088_));
 sky130_fd_sc_hd__a221o_1 _4162_ (.A1(\second_row[13][5] ),
    .A2(_1726_),
    .B1(_1907_),
    .B2(\second_row[5][5] ),
    .C1(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__a2111o_1 _4163_ (.A1(\second_row[1][5] ),
    .A2(_1938_),
    .B1(_2085_),
    .C1(_2087_),
    .D1(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__nor3_2 _4164_ (.A(_2083_),
    .B(_2084_),
    .C(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__o22ai_1 _4165_ (.A1(_2070_),
    .A2(_2080_),
    .B1(_2081_),
    .B2(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__nor2_1 _4166_ (.A(\second_row[0][4] ),
    .B(_1782_),
    .Y(_2093_));
 sky130_fd_sc_hd__a22o_1 _4167_ (.A1(\second_row[16][4] ),
    .A2(_1788_),
    .B1(_1804_),
    .B2(\second_row[8][4] ),
    .X(_2094_));
 sky130_fd_sc_hd__a221o_1 _4168_ (.A1(\second_row[9][4] ),
    .A2(_1799_),
    .B1(_1786_),
    .B2(\second_row[11][4] ),
    .C1(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__a221o_1 _4169_ (.A1(\second_row[15][4] ),
    .A2(_1933_),
    .B1(_1914_),
    .B2(\second_row[3][4] ),
    .C1(_1793_),
    .X(_2096_));
 sky130_fd_sc_hd__or2_1 _4170_ (.A(_2095_),
    .B(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__a22o_1 _4171_ (.A1(\second_row[1][4] ),
    .A2(_1936_),
    .B1(_1954_),
    .B2(\second_row[7][4] ),
    .X(_2098_));
 sky130_fd_sc_hd__a22o_1 _4172_ (.A1(\second_row[10][4] ),
    .A2(_1926_),
    .B1(_1791_),
    .B2(\second_row[17][4] ),
    .X(_2099_));
 sky130_fd_sc_hd__a221o_1 _4173_ (.A1(\second_row[5][4] ),
    .A2(_1906_),
    .B1(_1911_),
    .B2(\second_row[12][4] ),
    .C1(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__a22o_1 _4174_ (.A1(\second_row[6][4] ),
    .A2(_1829_),
    .B1(_1939_),
    .B2(\second_row[2][4] ),
    .X(_2101_));
 sky130_fd_sc_hd__a221o_1 _4175_ (.A1(\second_row[4][4] ),
    .A2(_1951_),
    .B1(_1923_),
    .B2(\second_row[14][4] ),
    .C1(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__a2111o_1 _4176_ (.A1(\second_row[13][4] ),
    .A2(_1726_),
    .B1(_2098_),
    .C1(_2100_),
    .D1(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__nor2_1 _4177_ (.A(_2097_),
    .B(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__a22o_1 _4178_ (.A1(\first_row[2][4] ),
    .A2(_1936_),
    .B1(_1829_),
    .B2(\first_row[7][4] ),
    .X(_2105_));
 sky130_fd_sc_hd__a221o_1 _4179_ (.A1(\first_row[15][4] ),
    .A2(_1923_),
    .B1(_1940_),
    .B2(\first_row[3][4] ),
    .C1(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__a22o_1 _4180_ (.A1(\first_row[17][4] ),
    .A2(_1943_),
    .B1(_1929_),
    .B2(\first_row[1][4] ),
    .X(_2107_));
 sky130_fd_sc_hd__a221o_1 _4181_ (.A1(\first_row[8][4] ),
    .A2(_1954_),
    .B1(_1927_),
    .B2(\first_row[11][4] ),
    .C1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__a2111o_1 _4182_ (.A1(\first_row[16][4] ),
    .A2(_1933_),
    .B1(_1919_),
    .C1(_2106_),
    .D1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__a22o_1 _4183_ (.A1(\first_row[13][4] ),
    .A2(_1911_),
    .B1(_1799_),
    .B2(\first_row[10][4] ),
    .X(_2110_));
 sky130_fd_sc_hd__a22o_1 _4184_ (.A1(\first_row[5][4] ),
    .A2(_1951_),
    .B1(_1914_),
    .B2(\first_row[4][4] ),
    .X(_2111_));
 sky130_fd_sc_hd__a22o_1 _4185_ (.A1(\first_row[14][4] ),
    .A2(_1726_),
    .B1(_1786_),
    .B2(\first_row[12][4] ),
    .X(_2112_));
 sky130_fd_sc_hd__a22o_1 _4186_ (.A1(\first_row[6][4] ),
    .A2(_1906_),
    .B1(_1804_),
    .B2(\first_row[9][4] ),
    .X(_2113_));
 sky130_fd_sc_hd__or4_2 _4187_ (.A(_2110_),
    .B(_2111_),
    .C(_2112_),
    .D(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__o22ai_2 _4188_ (.A1(\first_row[0][4] ),
    .A2(_1904_),
    .B1(_2109_),
    .B2(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__o21ai_1 _4189_ (.A1(_2093_),
    .A2(_2104_),
    .B1(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__nor2_1 _4190_ (.A(\first_row[0][3] ),
    .B(_1904_),
    .Y(_2117_));
 sky130_fd_sc_hd__a22o_1 _4191_ (.A1(\first_row[17][3] ),
    .A2(_1788_),
    .B1(_1785_),
    .B2(\first_row[12][3] ),
    .X(_2118_));
 sky130_fd_sc_hd__a221o_1 _4192_ (.A1(\first_row[4][3] ),
    .A2(_1914_),
    .B1(_1923_),
    .B2(\first_row[15][3] ),
    .C1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__a211o_1 _4193_ (.A1(\first_row[16][3] ),
    .A2(_1933_),
    .B1(_1919_),
    .C1(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__a22o_1 _4194_ (.A1(\first_row[6][3] ),
    .A2(_1826_),
    .B1(_1831_),
    .B2(\first_row[5][3] ),
    .X(_2121_));
 sky130_fd_sc_hd__a221o_1 _4195_ (.A1(\first_row[14][3] ),
    .A2(_1725_),
    .B1(_1954_),
    .B2(\first_row[8][3] ),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__a22o_1 _4196_ (.A1(\first_row[10][3] ),
    .A2(_1798_),
    .B1(_1817_),
    .B2(\first_row[11][3] ),
    .X(_2123_));
 sky130_fd_sc_hd__a221o_1 _4197_ (.A1(\first_row[9][3] ),
    .A2(_1804_),
    .B1(_1939_),
    .B2(\first_row[3][3] ),
    .C1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _4198_ (.A1(\first_row[13][3] ),
    .A2(_1819_),
    .B1(_1868_),
    .B2(\first_row[1][3] ),
    .X(_2125_));
 sky130_fd_sc_hd__a221o_1 _4199_ (.A1(\first_row[2][3] ),
    .A2(_1936_),
    .B1(_1829_),
    .B2(\first_row[7][3] ),
    .C1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__or3_1 _4200_ (.A(_2122_),
    .B(_2124_),
    .C(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__nor2_2 _4201_ (.A(_2120_),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__nor2_1 _4202_ (.A(\second_row[0][3] ),
    .B(_1782_),
    .Y(_2129_));
 sky130_fd_sc_hd__a22o_1 _4203_ (.A1(\second_row[13][3] ),
    .A2(_1726_),
    .B1(_1926_),
    .B2(\second_row[10][3] ),
    .X(_2130_));
 sky130_fd_sc_hd__a221o_1 _4204_ (.A1(\second_row[9][3] ),
    .A2(_1799_),
    .B1(_1786_),
    .B2(\second_row[11][3] ),
    .C1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__a221o_1 _4205_ (.A1(\second_row[5][3] ),
    .A2(_1906_),
    .B1(_1933_),
    .B2(\second_row[15][3] ),
    .C1(_1793_),
    .X(_2132_));
 sky130_fd_sc_hd__a22o_1 _4206_ (.A1(\second_row[7][3] ),
    .A2(_1954_),
    .B1(_1804_),
    .B2(\second_row[8][3] ),
    .X(_2133_));
 sky130_fd_sc_hd__a22o_1 _4207_ (.A1(\second_row[1][3] ),
    .A2(_1790_),
    .B1(_1791_),
    .B2(\second_row[17][3] ),
    .X(_2134_));
 sky130_fd_sc_hd__a221o_1 _4208_ (.A1(\second_row[16][3] ),
    .A2(_1788_),
    .B1(_1829_),
    .B2(\second_row[6][3] ),
    .C1(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__a22o_1 _4209_ (.A1(\second_row[12][3] ),
    .A2(_1819_),
    .B1(_1833_),
    .B2(\second_row[2][3] ),
    .X(_2136_));
 sky130_fd_sc_hd__a221o_1 _4210_ (.A1(\second_row[4][3] ),
    .A2(_1951_),
    .B1(_1923_),
    .B2(\second_row[14][3] ),
    .C1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__a2111o_1 _4211_ (.A1(\second_row[3][3] ),
    .A2(_1914_),
    .B1(_2133_),
    .C1(_2135_),
    .D1(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__nor3_2 _4212_ (.A(_2131_),
    .B(_2132_),
    .C(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__o22ai_4 _4213_ (.A1(_2117_),
    .A2(_2128_),
    .B1(_2129_),
    .B2(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__a22o_1 _4214_ (.A1(\second_row[7][1] ),
    .A2(_1813_),
    .B1(_1833_),
    .B2(\second_row[2][1] ),
    .X(_2141_));
 sky130_fd_sc_hd__a211o_1 _4215_ (.A1(\second_row[12][1] ),
    .A2(_1911_),
    .B1(_2141_),
    .C1(_1793_),
    .X(_2142_));
 sky130_fd_sc_hd__and3_1 _4216_ (.A(\second_row[9][1] ),
    .B(_1775_),
    .C(_1796_),
    .X(_2143_));
 sky130_fd_sc_hd__a221o_1 _4217_ (.A1(\second_row[16][1] ),
    .A2(_1788_),
    .B1(_1803_),
    .B2(\second_row[8][1] ),
    .C1(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__and3_1 _4218_ (.A(\second_row[14][1] ),
    .B(_1732_),
    .C(_1780_),
    .X(_2145_));
 sky130_fd_sc_hd__a221o_1 _4219_ (.A1(\second_row[13][1] ),
    .A2(_1725_),
    .B1(_1807_),
    .B2(\second_row[15][1] ),
    .C1(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__a22o_1 _4220_ (.A1(\second_row[5][1] ),
    .A2(_1826_),
    .B1(_1828_),
    .B2(\second_row[6][1] ),
    .X(_2147_));
 sky130_fd_sc_hd__a22o_1 _4221_ (.A1(\second_row[3][1] ),
    .A2(_1821_),
    .B1(_1785_),
    .B2(\second_row[11][1] ),
    .X(_2148_));
 sky130_fd_sc_hd__and3_1 _4222_ (.A(\second_row[1][1] ),
    .B(_1723_),
    .C(_1777_),
    .X(_2149_));
 sky130_fd_sc_hd__and3_1 _4223_ (.A(\second_row[17][1] ),
    .B(_1717_),
    .C(_1780_),
    .X(_2150_));
 sky130_fd_sc_hd__and3_1 _4224_ (.A(\second_row[4][1] ),
    .B(_1850_),
    .C(_1801_),
    .X(_2151_));
 sky130_fd_sc_hd__a2111o_1 _4225_ (.A1(\second_row[10][1] ),
    .A2(_1816_),
    .B1(_2149_),
    .C1(_2150_),
    .D1(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__or4_1 _4226_ (.A(_2146_),
    .B(_2147_),
    .C(_2148_),
    .D(_2152_),
    .X(_2153_));
 sky130_fd_sc_hd__o32a_2 _4227_ (.A1(_2142_),
    .A2(_2144_),
    .A3(_2153_),
    .B1(_1782_),
    .B2(\second_row[0][1] ),
    .X(_2154_));
 sky130_fd_sc_hd__a22o_1 _4228_ (.A1(\first_row[13][1] ),
    .A2(_1819_),
    .B1(_1868_),
    .B2(\first_row[1][1] ),
    .X(_2155_));
 sky130_fd_sc_hd__a221o_1 _4229_ (.A1(\first_row[2][1] ),
    .A2(_1790_),
    .B1(_1803_),
    .B2(\first_row[9][1] ),
    .C1(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__a21o_1 _4230_ (.A1(\first_row[16][1] ),
    .A2(_1808_),
    .B1(_1842_),
    .X(_2157_));
 sky130_fd_sc_hd__a22o_1 _4231_ (.A1(\first_row[11][1] ),
    .A2(_1817_),
    .B1(_1833_),
    .B2(\first_row[3][1] ),
    .X(_2158_));
 sky130_fd_sc_hd__a22o_1 _4232_ (.A1(\first_row[5][1] ),
    .A2(_1831_),
    .B1(_1810_),
    .B2(\first_row[15][1] ),
    .X(_2159_));
 sky130_fd_sc_hd__and3_1 _4233_ (.A(\first_row[6][1] ),
    .B(_1723_),
    .C(_1820_),
    .X(_2160_));
 sky130_fd_sc_hd__and3_1 _4234_ (.A(\first_row[14][1] ),
    .B(_1718_),
    .C(_1723_),
    .X(_2161_));
 sky130_fd_sc_hd__and3_1 _4235_ (.A(\first_row[10][1] ),
    .B(_1775_),
    .C(_1796_),
    .X(_2162_));
 sky130_fd_sc_hd__a2111o_1 _4236_ (.A1(\first_row[17][1] ),
    .A2(_1787_),
    .B1(_2160_),
    .C1(_2161_),
    .D1(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__and3_1 _4237_ (.A(\first_row[12][1] ),
    .B(_1718_),
    .C(_1853_),
    .X(_2164_));
 sky130_fd_sc_hd__and3_1 _4238_ (.A(\first_row[4][1] ),
    .B(_1850_),
    .C(_1853_),
    .X(_2165_));
 sky130_fd_sc_hd__and3_1 _4239_ (.A(\first_row[8][1] ),
    .B(_1853_),
    .C(_1796_),
    .X(_2166_));
 sky130_fd_sc_hd__a2111o_1 _4240_ (.A1(\first_row[7][1] ),
    .A2(_1828_),
    .B1(_2164_),
    .C1(_2165_),
    .D1(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__or4_2 _4241_ (.A(_2158_),
    .B(_2159_),
    .C(_2163_),
    .D(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__o32a_1 _4242_ (.A1(_2156_),
    .A2(_2157_),
    .A3(_2168_),
    .B1(_1857_),
    .B2(\first_row[0][1] ),
    .X(_2169_));
 sky130_fd_sc_hd__xor2_2 _4243_ (.A(_2154_),
    .B(_2169_),
    .X(_2170_));
 sky130_fd_sc_hd__a32o_1 _4244_ (.A1(_1860_),
    .A2(_1858_),
    .A3(_2170_),
    .B1(_2169_),
    .B2(_2154_),
    .X(_2171_));
 sky130_fd_sc_hd__a22o_1 _4245_ (.A1(\first_row[17][2] ),
    .A2(_1788_),
    .B1(_1828_),
    .B2(\first_row[7][2] ),
    .X(_2172_));
 sky130_fd_sc_hd__a221o_1 _4246_ (.A1(\first_row[2][2] ),
    .A2(_1790_),
    .B1(_1926_),
    .B2(\first_row[11][2] ),
    .C1(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__a22o_1 _4247_ (.A1(\first_row[15][2] ),
    .A2(_1810_),
    .B1(_1868_),
    .B2(\first_row[1][2] ),
    .X(_2174_));
 sky130_fd_sc_hd__a221o_1 _4248_ (.A1(\first_row[8][2] ),
    .A2(_1954_),
    .B1(_1939_),
    .B2(\first_row[3][2] ),
    .C1(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__a2111o_1 _4249_ (.A1(\first_row[16][2] ),
    .A2(_1808_),
    .B1(_1842_),
    .C1(_2173_),
    .D1(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__a22o_1 _4250_ (.A1(\first_row[13][2] ),
    .A2(_1819_),
    .B1(_1822_),
    .B2(\first_row[4][2] ),
    .X(_2177_));
 sky130_fd_sc_hd__a221o_1 _4251_ (.A1(\first_row[12][2] ),
    .A2(_1786_),
    .B1(_1804_),
    .B2(\first_row[9][2] ),
    .C1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__a22o_1 _4252_ (.A1(\first_row[6][2] ),
    .A2(_1826_),
    .B1(_1798_),
    .B2(\first_row[10][2] ),
    .X(_2179_));
 sky130_fd_sc_hd__a221o_1 _4253_ (.A1(\first_row[14][2] ),
    .A2(_1725_),
    .B1(_1951_),
    .B2(\first_row[5][2] ),
    .C1(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__or2_1 _4254_ (.A(_2178_),
    .B(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__o22a_1 _4255_ (.A1(\first_row[0][2] ),
    .A2(_1904_),
    .B1(_2176_),
    .B2(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__a22o_1 _4256_ (.A1(\second_row[5][2] ),
    .A2(_1906_),
    .B1(_1803_),
    .B2(\second_row[8][2] ),
    .X(_2183_));
 sky130_fd_sc_hd__a221o_1 _4257_ (.A1(\second_row[10][2] ),
    .A2(_1926_),
    .B1(_1786_),
    .B2(\second_row[11][2] ),
    .C1(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__a22o_1 _4258_ (.A1(\second_row[1][2] ),
    .A2(_1936_),
    .B1(_1788_),
    .B2(\second_row[16][2] ),
    .X(_2185_));
 sky130_fd_sc_hd__a22o_1 _4259_ (.A1(\second_row[15][2] ),
    .A2(_1808_),
    .B1(_1923_),
    .B2(\second_row[14][2] ),
    .X(_2186_));
 sky130_fd_sc_hd__a211o_1 _4260_ (.A1(\second_row[17][2] ),
    .A2(_1791_),
    .B1(_2185_),
    .C1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__a22o_1 _4261_ (.A1(\second_row[9][2] ),
    .A2(_1798_),
    .B1(_1833_),
    .B2(\second_row[2][2] ),
    .X(_2188_));
 sky130_fd_sc_hd__a221o_1 _4262_ (.A1(\second_row[4][2] ),
    .A2(_1831_),
    .B1(_1911_),
    .B2(\second_row[12][2] ),
    .C1(_2188_),
    .X(_2189_));
 sky130_fd_sc_hd__a22o_1 _4263_ (.A1(\second_row[7][2] ),
    .A2(_1813_),
    .B1(_1828_),
    .B2(\second_row[6][2] ),
    .X(_2190_));
 sky130_fd_sc_hd__a221o_1 _4264_ (.A1(\second_row[13][2] ),
    .A2(_1725_),
    .B1(_1822_),
    .B2(\second_row[3][2] ),
    .C1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__or3_1 _4265_ (.A(_1793_),
    .B(_2189_),
    .C(_2191_),
    .X(_2192_));
 sky130_fd_sc_hd__o32a_2 _4266_ (.A1(_2184_),
    .A2(_2187_),
    .A3(_2192_),
    .B1(_1782_),
    .B2(\second_row[0][2] ),
    .X(_2193_));
 sky130_fd_sc_hd__xor2_2 _4267_ (.A(_2182_),
    .B(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__nor4_1 _4268_ (.A(_2117_),
    .B(_2128_),
    .C(_2129_),
    .D(_2139_),
    .Y(_2195_));
 sky130_fd_sc_hd__and2_1 _4269_ (.A(_2182_),
    .B(_2193_),
    .X(_2196_));
 sky130_fd_sc_hd__a211o_1 _4270_ (.A1(_2171_),
    .A2(_2194_),
    .B1(_2195_),
    .C1(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__nor2_1 _4271_ (.A(_2093_),
    .B(_2104_),
    .Y(_2198_));
 sky130_fd_sc_hd__and2b_1 _4272_ (.A_N(_2115_),
    .B(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__a31o_1 _4273_ (.A1(_2116_),
    .A2(_2140_),
    .A3(_2197_),
    .B1(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__nor4_1 _4274_ (.A(_2070_),
    .B(_2080_),
    .C(_2081_),
    .D(_2091_),
    .Y(_2201_));
 sky130_fd_sc_hd__a21o_1 _4275_ (.A1(_2092_),
    .A2(_2200_),
    .B1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__nor2_1 _4276_ (.A(\first_row[0][6] ),
    .B(_1904_),
    .Y(_2203_));
 sky130_fd_sc_hd__a22o_1 _4277_ (.A1(\first_row[10][6] ),
    .A2(_1945_),
    .B1(_1909_),
    .B2(\first_row[9][6] ),
    .X(_2204_));
 sky130_fd_sc_hd__a221o_1 _4278_ (.A1(\first_row[14][6] ),
    .A2(_1727_),
    .B1(_1956_),
    .B2(\first_row[8][6] ),
    .C1(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__a22o_1 _4279_ (.A1(\first_row[2][6] ),
    .A2(_1937_),
    .B1(_1943_),
    .B2(\first_row[17][6] ),
    .X(_2206_));
 sky130_fd_sc_hd__a221o_1 _4280_ (.A1(\first_row[11][6] ),
    .A2(_1927_),
    .B1(_1922_),
    .B2(\first_row[7][6] ),
    .C1(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__a22o_1 _4281_ (.A1(\first_row[15][6] ),
    .A2(_1924_),
    .B1(_1929_),
    .B2(\first_row[1][6] ),
    .X(_2208_));
 sky130_fd_sc_hd__a221o_1 _4282_ (.A1(\first_row[12][6] ),
    .A2(_1949_),
    .B1(_1940_),
    .B2(\first_row[3][6] ),
    .C1(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__a2111o_1 _4283_ (.A1(\first_row[16][6] ),
    .A2(_1934_),
    .B1(_1920_),
    .C1(_2207_),
    .D1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _4284_ (.A1(\first_row[6][6] ),
    .A2(_1907_),
    .B1(_1912_),
    .B2(\first_row[13][6] ),
    .X(_2211_));
 sky130_fd_sc_hd__a221o_1 _4285_ (.A1(\first_row[5][6] ),
    .A2(_1953_),
    .B1(_1916_),
    .B2(\first_row[4][6] ),
    .C1(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__nor3_1 _4286_ (.A(_2205_),
    .B(_2210_),
    .C(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__nor2_1 _4287_ (.A(\second_row[0][6] ),
    .B(_1782_),
    .Y(_2214_));
 sky130_fd_sc_hd__a22o_1 _4288_ (.A1(\second_row[4][6] ),
    .A2(_1952_),
    .B1(_1924_),
    .B2(\second_row[14][6] ),
    .X(_2215_));
 sky130_fd_sc_hd__a221o_1 _4289_ (.A1(\second_row[5][6] ),
    .A2(_1908_),
    .B1(_1913_),
    .B2(\second_row[12][6] ),
    .C1(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__a221o_1 _4290_ (.A1(\second_row[15][6] ),
    .A2(_1934_),
    .B1(_1928_),
    .B2(\second_row[10][6] ),
    .C1(_1793_),
    .X(_2217_));
 sky130_fd_sc_hd__a22o_1 _4291_ (.A1(\second_row[13][6] ),
    .A2(_1727_),
    .B1(_1949_),
    .B2(\second_row[11][6] ),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_1 _4292_ (.A1(\second_row[3][6] ),
    .A2(_1915_),
    .B1(_1791_),
    .B2(\second_row[17][6] ),
    .X(_2219_));
 sky130_fd_sc_hd__a221o_1 _4293_ (.A1(\second_row[1][6] ),
    .A2(_1937_),
    .B1(_1943_),
    .B2(\second_row[16][6] ),
    .C1(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__a22o_1 _4294_ (.A1(\second_row[9][6] ),
    .A2(_1945_),
    .B1(_1921_),
    .B2(\second_row[6][6] ),
    .X(_2221_));
 sky130_fd_sc_hd__a221o_1 _4295_ (.A1(\second_row[7][6] ),
    .A2(_1955_),
    .B1(_1940_),
    .B2(\second_row[2][6] ),
    .C1(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__a2111o_1 _4296_ (.A1(\second_row[8][6] ),
    .A2(_1910_),
    .B1(_2218_),
    .C1(_2220_),
    .D1(_2222_),
    .X(_2223_));
 sky130_fd_sc_hd__nor3_1 _4297_ (.A(_2216_),
    .B(_2217_),
    .C(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__o22ai_1 _4298_ (.A1(_2203_),
    .A2(_2213_),
    .B1(_2214_),
    .B2(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nor4_1 _4299_ (.A(_2203_),
    .B(_2213_),
    .C(_2214_),
    .D(_2224_),
    .Y(_2226_));
 sky130_fd_sc_hd__a21o_1 _4300_ (.A1(_2202_),
    .A2(_2225_),
    .B1(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__nor2_1 _4301_ (.A(_2069_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__nor2_1 _4302_ (.A(\second_row[0][7] ),
    .B(_1865_),
    .Y(_2229_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(\second_row[3][7] ),
    .A2(_1938_),
    .B1(_1941_),
    .B2(\second_row[4][7] ),
    .X(_2230_));
 sky130_fd_sc_hd__a22o_1 _4304_ (.A1(\second_row[7][7] ),
    .A2(_1908_),
    .B1(_1877_),
    .B2(\second_row[1][7] ),
    .X(_2231_));
 sky130_fd_sc_hd__a221o_1 _4305_ (.A1(\second_row[14][7] ),
    .A2(_1913_),
    .B1(_1922_),
    .B2(\second_row[8][7] ),
    .C1(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__a22o_1 _4306_ (.A1(\second_row[11][7] ),
    .A2(_1945_),
    .B1(_1909_),
    .B2(\second_row[10][7] ),
    .X(_2233_));
 sky130_fd_sc_hd__a221o_1 _4307_ (.A1(\second_row[6][7] ),
    .A2(_1952_),
    .B1(_1915_),
    .B2(\second_row[5][7] ),
    .C1(_2233_),
    .X(_2234_));
 sky130_fd_sc_hd__a22o_1 _4308_ (.A1(\second_row[15][7] ),
    .A2(_1727_),
    .B1(_1925_),
    .B2(\second_row[16][7] ),
    .X(_2235_));
 sky130_fd_sc_hd__a221o_1 _4309_ (.A1(\second_row[9][7] ),
    .A2(_1955_),
    .B1(_1928_),
    .B2(\second_row[12][7] ),
    .C1(_1866_),
    .X(_2236_));
 sky130_fd_sc_hd__a2111o_1 _4310_ (.A1(\second_row[17][7] ),
    .A2(_1935_),
    .B1(_2234_),
    .C1(_2235_),
    .D1(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__a211o_1 _4311_ (.A1(\second_row[13][7] ),
    .A2(_1950_),
    .B1(_2232_),
    .C1(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__a211oi_2 _4312_ (.A1(\second_row[2][7] ),
    .A2(_1930_),
    .B1(_2230_),
    .C1(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__a22o_1 _4313_ (.A1(\third_row[4][7] ),
    .A2(_1915_),
    .B1(_1949_),
    .B2(\third_row[12][7] ),
    .X(_2240_));
 sky130_fd_sc_hd__a221o_1 _4314_ (.A1(\third_row[8][7] ),
    .A2(_1956_),
    .B1(_1946_),
    .B2(\third_row[10][7] ),
    .C1(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__a22o_1 _4315_ (.A1(\third_row[13][7] ),
    .A2(_1912_),
    .B1(_1909_),
    .B2(\third_row[9][7] ),
    .X(_2242_));
 sky130_fd_sc_hd__a221o_1 _4316_ (.A1(\third_row[14][7] ),
    .A2(_1728_),
    .B1(_1953_),
    .B2(\third_row[5][7] ),
    .C1(_2242_),
    .X(_2243_));
 sky130_fd_sc_hd__a22o_1 _4317_ (.A1(\third_row[2][7] ),
    .A2(_1937_),
    .B1(_1940_),
    .B2(\third_row[3][7] ),
    .X(_2244_));
 sky130_fd_sc_hd__a221o_1 _4318_ (.A1(\third_row[6][7] ),
    .A2(_1907_),
    .B1(_1944_),
    .B2(\third_row[17][7] ),
    .C1(_2244_),
    .X(_2245_));
 sky130_fd_sc_hd__a22o_1 _4319_ (.A1(\third_row[7][7] ),
    .A2(_1921_),
    .B1(_1924_),
    .B2(\third_row[15][7] ),
    .X(_2246_));
 sky130_fd_sc_hd__a221o_1 _4320_ (.A1(\third_row[11][7] ),
    .A2(_1927_),
    .B1(_1930_),
    .B2(\third_row[1][7] ),
    .C1(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__a2111o_1 _4321_ (.A1(\third_row[16][7] ),
    .A2(_1935_),
    .B1(_1920_),
    .C1(_2245_),
    .D1(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__or3_1 _4322_ (.A(_2241_),
    .B(_2243_),
    .C(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__o21ai_1 _4323_ (.A1(\third_row[0][7] ),
    .A2(_1905_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__o21a_1 _4324_ (.A1(_2229_),
    .A2(_2239_),
    .B1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__nor3_1 _4325_ (.A(_2250_),
    .B(_2229_),
    .C(_2239_),
    .Y(_2252_));
 sky130_fd_sc_hd__nor2_1 _4326_ (.A(\third_row[0][5] ),
    .B(_1904_),
    .Y(_2253_));
 sky130_fd_sc_hd__a22o_1 _4327_ (.A1(\third_row[12][5] ),
    .A2(_1949_),
    .B1(_1909_),
    .B2(\third_row[9][5] ),
    .X(_2254_));
 sky130_fd_sc_hd__a221o_1 _4328_ (.A1(\third_row[13][5] ),
    .A2(_1912_),
    .B1(_1916_),
    .B2(\third_row[4][5] ),
    .C1(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__a22o_1 _4329_ (.A1(\third_row[17][5] ),
    .A2(_1943_),
    .B1(_1940_),
    .B2(\third_row[3][5] ),
    .X(_2256_));
 sky130_fd_sc_hd__a221o_1 _4330_ (.A1(\third_row[11][5] ),
    .A2(_1927_),
    .B1(_1929_),
    .B2(\third_row[1][5] ),
    .C1(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__a22o_1 _4331_ (.A1(\third_row[2][5] ),
    .A2(_1937_),
    .B1(_1921_),
    .B2(\third_row[7][5] ),
    .X(_2258_));
 sky130_fd_sc_hd__a221o_1 _4332_ (.A1(\third_row[10][5] ),
    .A2(_1945_),
    .B1(_1924_),
    .B2(\third_row[15][5] ),
    .C1(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__a2111o_1 _4333_ (.A1(\third_row[16][5] ),
    .A2(_1934_),
    .B1(_1919_),
    .C1(_2257_),
    .D1(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a22o_1 _4334_ (.A1(\third_row[6][5] ),
    .A2(_1907_),
    .B1(_1955_),
    .B2(\third_row[8][5] ),
    .X(_2261_));
 sky130_fd_sc_hd__a221o_1 _4335_ (.A1(\third_row[14][5] ),
    .A2(_1727_),
    .B1(_1952_),
    .B2(\third_row[5][5] ),
    .C1(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__nor3_2 _4336_ (.A(_2255_),
    .B(_2260_),
    .C(_2262_),
    .Y(_2263_));
 sky130_fd_sc_hd__a221o_1 _4337_ (.A1(\second_row[15][5] ),
    .A2(_1727_),
    .B1(_1934_),
    .B2(\second_row[17][5] ),
    .C1(_1866_),
    .X(_2264_));
 sky130_fd_sc_hd__a22o_1 _4338_ (.A1(\second_row[11][5] ),
    .A2(_1799_),
    .B1(_1929_),
    .B2(\second_row[2][5] ),
    .X(_2265_));
 sky130_fd_sc_hd__a221o_1 _4339_ (.A1(\second_row[9][5] ),
    .A2(_1955_),
    .B1(_1924_),
    .B2(\second_row[16][5] ),
    .C1(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__and3_1 _4340_ (.A(\second_row[8][5] ),
    .B(_1796_),
    .C(_1815_),
    .X(_2267_));
 sky130_fd_sc_hd__a221o_1 _4341_ (.A1(\second_row[3][5] ),
    .A2(_1937_),
    .B1(_1949_),
    .B2(\second_row[13][5] ),
    .C1(_2267_),
    .X(_2268_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(\second_row[6][5] ),
    .A2(_1951_),
    .B1(_1804_),
    .B2(\second_row[10][5] ),
    .X(_2269_));
 sky130_fd_sc_hd__a221o_1 _4343_ (.A1(\second_row[7][5] ),
    .A2(_1906_),
    .B1(_1912_),
    .B2(\second_row[14][5] ),
    .C1(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(\second_row[4][5] ),
    .A2(_1939_),
    .B1(_1877_),
    .B2(\second_row[1][5] ),
    .X(_2271_));
 sky130_fd_sc_hd__a221o_1 _4345_ (.A1(\second_row[12][5] ),
    .A2(_1927_),
    .B1(_1915_),
    .B2(\second_row[5][5] ),
    .C1(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__or4_2 _4346_ (.A(_2266_),
    .B(_2268_),
    .C(_2270_),
    .D(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__o22ai_1 _4347_ (.A1(\second_row[0][5] ),
    .A2(_1865_),
    .B1(_2264_),
    .B2(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__o21ai_1 _4348_ (.A1(_2253_),
    .A2(_2263_),
    .B1(_2274_),
    .Y(_2275_));
 sky130_fd_sc_hd__nor2_1 _4349_ (.A(\third_row[0][4] ),
    .B(_1904_),
    .Y(_2276_));
 sky130_fd_sc_hd__a22o_1 _4350_ (.A1(\third_row[8][4] ),
    .A2(_1954_),
    .B1(_1786_),
    .B2(\third_row[12][4] ),
    .X(_2277_));
 sky130_fd_sc_hd__a221o_1 _4351_ (.A1(\third_row[5][4] ),
    .A2(_1952_),
    .B1(_1804_),
    .B2(\third_row[9][4] ),
    .C1(_2277_),
    .X(_2278_));
 sky130_fd_sc_hd__a22o_1 _4352_ (.A1(\third_row[15][4] ),
    .A2(_1923_),
    .B1(_1868_),
    .B2(\third_row[1][4] ),
    .X(_2279_));
 sky130_fd_sc_hd__a221o_1 _4353_ (.A1(\third_row[11][4] ),
    .A2(_1926_),
    .B1(_1829_),
    .B2(\third_row[7][4] ),
    .C1(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__a22o_1 _4354_ (.A1(\third_row[17][4] ),
    .A2(_1788_),
    .B1(_1799_),
    .B2(\third_row[10][4] ),
    .X(_2281_));
 sky130_fd_sc_hd__a221o_1 _4355_ (.A1(\third_row[2][4] ),
    .A2(_1936_),
    .B1(_1939_),
    .B2(\third_row[3][4] ),
    .C1(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__a2111o_1 _4356_ (.A1(\third_row[16][4] ),
    .A2(_1933_),
    .B1(_1919_),
    .C1(_2280_),
    .D1(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__a22o_1 _4357_ (.A1(\third_row[13][4] ),
    .A2(_1911_),
    .B1(_1914_),
    .B2(\third_row[4][4] ),
    .X(_2284_));
 sky130_fd_sc_hd__a221o_1 _4358_ (.A1(\third_row[14][4] ),
    .A2(_1726_),
    .B1(_1907_),
    .B2(\third_row[6][4] ),
    .C1(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__nor3_2 _4359_ (.A(_2278_),
    .B(_2283_),
    .C(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__a221o_1 _4360_ (.A1(\second_row[15][4] ),
    .A2(_1726_),
    .B1(_1933_),
    .B2(\second_row[17][4] ),
    .C1(_1866_),
    .X(_2287_));
 sky130_fd_sc_hd__a22o_1 _4361_ (.A1(\second_row[3][4] ),
    .A2(_1936_),
    .B1(_1951_),
    .B2(\second_row[6][4] ),
    .X(_2288_));
 sky130_fd_sc_hd__a221o_1 _4362_ (.A1(\second_row[7][4] ),
    .A2(_1906_),
    .B1(_1829_),
    .B2(\second_row[8][4] ),
    .C1(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__and3_1 _4363_ (.A(\second_row[13][4] ),
    .B(_1719_),
    .C(_1853_),
    .X(_2290_));
 sky130_fd_sc_hd__a221o_1 _4364_ (.A1(\second_row[9][4] ),
    .A2(_1954_),
    .B1(_1929_),
    .B2(\second_row[2][4] ),
    .C1(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__a22o_1 _4365_ (.A1(\second_row[11][4] ),
    .A2(_1799_),
    .B1(_1939_),
    .B2(\second_row[4][4] ),
    .X(_2292_));
 sky130_fd_sc_hd__a221o_1 _4366_ (.A1(\second_row[14][4] ),
    .A2(_1911_),
    .B1(_1926_),
    .B2(\second_row[12][4] ),
    .C1(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__a22o_1 _4367_ (.A1(\second_row[5][4] ),
    .A2(_1914_),
    .B1(_1877_),
    .B2(\second_row[1][4] ),
    .X(_2294_));
 sky130_fd_sc_hd__a221o_1 _4368_ (.A1(\second_row[16][4] ),
    .A2(_1923_),
    .B1(_1804_),
    .B2(\second_row[10][4] ),
    .C1(_2294_),
    .X(_2295_));
 sky130_fd_sc_hd__or4_2 _4369_ (.A(_2289_),
    .B(_2291_),
    .C(_2293_),
    .D(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__o22ai_2 _4370_ (.A1(\second_row[0][4] ),
    .A2(_1865_),
    .B1(_2287_),
    .B2(_2296_),
    .Y(_2297_));
 sky130_fd_sc_hd__o21ai_2 _4371_ (.A1(_2276_),
    .A2(_2286_),
    .B1(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__and3_1 _4372_ (.A(\third_row[1][1] ),
    .B(_1777_),
    .C(_1801_),
    .X(_2299_));
 sky130_fd_sc_hd__and3_1 _4373_ (.A(\third_row[7][1] ),
    .B(_1796_),
    .C(_1815_),
    .X(_2300_));
 sky130_fd_sc_hd__and3_1 _4374_ (.A(\third_row[11][1] ),
    .B(_1719_),
    .C(_1815_),
    .X(_2301_));
 sky130_fd_sc_hd__a2111o_1 _4375_ (.A1(\third_row[17][1] ),
    .A2(_1787_),
    .B1(_2299_),
    .C1(_2300_),
    .D1(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__and3_1 _4376_ (.A(\third_row[3][1] ),
    .B(_1850_),
    .C(_1815_),
    .X(_2303_));
 sky130_fd_sc_hd__and3_1 _4377_ (.A(\third_row[14][1] ),
    .B(_1719_),
    .C(_1775_),
    .X(_2304_));
 sky130_fd_sc_hd__and3_1 _4378_ (.A(\third_row[2][1] ),
    .B(_1775_),
    .C(_1777_),
    .X(_2305_));
 sky130_fd_sc_hd__a2111o_1 _4379_ (.A1(\third_row[15][1] ),
    .A2(_1810_),
    .B1(_2303_),
    .C1(_2304_),
    .D1(_2305_),
    .X(_2306_));
 sky130_fd_sc_hd__a2111o_1 _4380_ (.A1(\third_row[16][1] ),
    .A2(_1807_),
    .B1(_1842_),
    .C1(_2302_),
    .D1(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__a22o_1 _4381_ (.A1(\third_row[10][1] ),
    .A2(_1798_),
    .B1(_1822_),
    .B2(\third_row[4][1] ),
    .X(_2308_));
 sky130_fd_sc_hd__a221o_1 _4382_ (.A1(\third_row[5][1] ),
    .A2(_1831_),
    .B1(_1785_),
    .B2(\third_row[12][1] ),
    .C1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__a22o_1 _4383_ (.A1(\third_row[6][1] ),
    .A2(_1826_),
    .B1(_1802_),
    .B2(\third_row[9][1] ),
    .X(_2310_));
 sky130_fd_sc_hd__a221o_1 _4384_ (.A1(\third_row[8][1] ),
    .A2(_1813_),
    .B1(_1819_),
    .B2(\third_row[13][1] ),
    .C1(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__o32a_4 _4385_ (.A1(_2307_),
    .A2(_2309_),
    .A3(_2311_),
    .B1(_1857_),
    .B2(\third_row[0][1] ),
    .X(_2312_));
 sky130_fd_sc_hd__a22o_1 _4386_ (.A1(\second_row[7][1] ),
    .A2(_1826_),
    .B1(_1813_),
    .B2(\second_row[9][1] ),
    .X(_2313_));
 sky130_fd_sc_hd__a22o_1 _4387_ (.A1(\second_row[13][1] ),
    .A2(_1785_),
    .B1(_1802_),
    .B2(\second_row[10][1] ),
    .X(_2314_));
 sky130_fd_sc_hd__a22o_1 _4388_ (.A1(\second_row[12][1] ),
    .A2(_1817_),
    .B1(_1822_),
    .B2(\second_row[5][1] ),
    .X(_2315_));
 sky130_fd_sc_hd__or4_1 _4389_ (.A(_1866_),
    .B(_2313_),
    .C(_2314_),
    .D(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(\second_row[15][1] ),
    .B(_1719_),
    .C(_1775_),
    .X(_2317_));
 sky130_fd_sc_hd__a221o_1 _4391_ (.A1(\second_row[17][1] ),
    .A2(_1807_),
    .B1(_1810_),
    .B2(\second_row[16][1] ),
    .C1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__a22o_1 _4392_ (.A1(\second_row[3][1] ),
    .A2(_1790_),
    .B1(_1828_),
    .B2(\second_row[8][1] ),
    .X(_2319_));
 sky130_fd_sc_hd__a22o_1 _4393_ (.A1(\second_row[6][1] ),
    .A2(_1831_),
    .B1(_1867_),
    .B2(\second_row[2][1] ),
    .X(_2320_));
 sky130_fd_sc_hd__and3_1 _4394_ (.A(\second_row[4][1] ),
    .B(_1850_),
    .C(_1815_),
    .X(_2321_));
 sky130_fd_sc_hd__and3_1 _4395_ (.A(\second_row[14][1] ),
    .B(_1719_),
    .C(_1801_),
    .X(_2322_));
 sky130_fd_sc_hd__and3_1 _4396_ (.A(\second_row[1][1] ),
    .B(_1777_),
    .C(_1853_),
    .X(_2323_));
 sky130_fd_sc_hd__a2111o_1 _4397_ (.A1(\second_row[11][1] ),
    .A2(_1797_),
    .B1(_2321_),
    .C1(_2322_),
    .D1(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__or4_1 _4398_ (.A(_2318_),
    .B(_2319_),
    .C(_2320_),
    .D(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__o22a_2 _4399_ (.A1(\second_row[0][1] ),
    .A2(_1865_),
    .B1(_2316_),
    .B2(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__xor2_2 _4400_ (.A(_2312_),
    .B(_2326_),
    .X(_2327_));
 sky130_fd_sc_hd__a32o_1 _4401_ (.A1(_1896_),
    .A2(_1898_),
    .A3(_2327_),
    .B1(_2326_),
    .B2(_2312_),
    .X(_2328_));
 sky130_fd_sc_hd__a22o_1 _4402_ (.A1(\third_row[13][2] ),
    .A2(_1819_),
    .B1(_1785_),
    .B2(\third_row[12][2] ),
    .X(_2329_));
 sky130_fd_sc_hd__a221o_1 _4403_ (.A1(\third_row[4][2] ),
    .A2(_1822_),
    .B1(_1833_),
    .B2(\third_row[3][2] ),
    .C1(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__a211o_1 _4404_ (.A1(\third_row[16][2] ),
    .A2(_1808_),
    .B1(_1919_),
    .C1(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__a22o_1 _4405_ (.A1(\third_row[8][2] ),
    .A2(_1813_),
    .B1(_1817_),
    .B2(\third_row[11][2] ),
    .X(_2332_));
 sky130_fd_sc_hd__a221o_1 _4406_ (.A1(\third_row[2][2] ),
    .A2(_1790_),
    .B1(_1798_),
    .B2(\third_row[10][2] ),
    .C1(_2332_),
    .X(_2333_));
 sky130_fd_sc_hd__a22o_1 _4407_ (.A1(\third_row[6][2] ),
    .A2(_1826_),
    .B1(_1828_),
    .B2(\third_row[7][2] ),
    .X(_2334_));
 sky130_fd_sc_hd__a221o_1 _4408_ (.A1(\third_row[17][2] ),
    .A2(_1788_),
    .B1(_1803_),
    .B2(\third_row[9][2] ),
    .C1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__a22o_1 _4409_ (.A1(\third_row[14][2] ),
    .A2(_1725_),
    .B1(_1810_),
    .B2(\third_row[15][2] ),
    .X(_2336_));
 sky130_fd_sc_hd__a221o_1 _4410_ (.A1(\third_row[5][2] ),
    .A2(_1951_),
    .B1(_1868_),
    .B2(\third_row[1][2] ),
    .C1(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__or3_2 _4411_ (.A(_2333_),
    .B(_2335_),
    .C(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__o22a_1 _4412_ (.A1(\third_row[0][2] ),
    .A2(_1857_),
    .B1(_2331_),
    .B2(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__a221o_1 _4413_ (.A1(\second_row[15][2] ),
    .A2(_1726_),
    .B1(_1808_),
    .B2(\second_row[17][2] ),
    .C1(_1866_),
    .X(_2340_));
 sky130_fd_sc_hd__a22o_1 _4414_ (.A1(\second_row[14][2] ),
    .A2(_1818_),
    .B1(_1868_),
    .B2(\second_row[2][2] ),
    .X(_2341_));
 sky130_fd_sc_hd__a221o_1 _4415_ (.A1(\second_row[7][2] ),
    .A2(_1826_),
    .B1(_1817_),
    .B2(\second_row[12][2] ),
    .C1(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__a22o_1 _4416_ (.A1(\second_row[9][2] ),
    .A2(_1813_),
    .B1(_1828_),
    .B2(\second_row[8][2] ),
    .X(_2343_));
 sky130_fd_sc_hd__a221o_1 _4417_ (.A1(\second_row[5][2] ),
    .A2(_1822_),
    .B1(_1803_),
    .B2(\second_row[10][2] ),
    .C1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__and3_1 _4418_ (.A(\second_row[1][2] ),
    .B(_1777_),
    .C(_1853_),
    .X(_2345_));
 sky130_fd_sc_hd__a221o_1 _4419_ (.A1(\second_row[3][2] ),
    .A2(_1790_),
    .B1(_1833_),
    .B2(\second_row[4][2] ),
    .C1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__a22o_1 _4420_ (.A1(\second_row[6][2] ),
    .A2(_1831_),
    .B1(_1785_),
    .B2(\second_row[13][2] ),
    .X(_2347_));
 sky130_fd_sc_hd__a221o_1 _4421_ (.A1(\second_row[11][2] ),
    .A2(_1798_),
    .B1(_1810_),
    .B2(\second_row[16][2] ),
    .C1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__or4_1 _4422_ (.A(_2342_),
    .B(_2344_),
    .C(_2346_),
    .D(_2348_),
    .X(_2349_));
 sky130_fd_sc_hd__o22a_1 _4423_ (.A1(\second_row[0][2] ),
    .A2(_1865_),
    .B1(_2340_),
    .B2(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__xor2_1 _4424_ (.A(_2339_),
    .B(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__nand2_1 _4425_ (.A(_2339_),
    .B(_2350_),
    .Y(_2352_));
 sky130_fd_sc_hd__a21bo_1 _4426_ (.A1(_2328_),
    .A2(_2351_),
    .B1_N(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__a22o_1 _4427_ (.A1(\third_row[8][3] ),
    .A2(_1954_),
    .B1(_1926_),
    .B2(\third_row[11][3] ),
    .X(_2354_));
 sky130_fd_sc_hd__a221o_1 _4428_ (.A1(\third_row[17][3] ),
    .A2(_1943_),
    .B1(_1911_),
    .B2(\third_row[13][3] ),
    .C1(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__a211o_1 _4429_ (.A1(\third_row[16][3] ),
    .A2(_1933_),
    .B1(_1919_),
    .C1(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__a22o_1 _4430_ (.A1(\third_row[6][3] ),
    .A2(_1906_),
    .B1(_1810_),
    .B2(\third_row[15][3] ),
    .X(_2357_));
 sky130_fd_sc_hd__a221o_1 _4431_ (.A1(\third_row[7][3] ),
    .A2(_1829_),
    .B1(_1868_),
    .B2(\third_row[1][3] ),
    .C1(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__a22o_1 _4432_ (.A1(\third_row[14][3] ),
    .A2(_1725_),
    .B1(_1803_),
    .B2(\third_row[9][3] ),
    .X(_2359_));
 sky130_fd_sc_hd__a221o_1 _4433_ (.A1(\third_row[2][3] ),
    .A2(_1936_),
    .B1(_1914_),
    .B2(\third_row[4][3] ),
    .C1(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__a22o_1 _4434_ (.A1(\third_row[10][3] ),
    .A2(_1799_),
    .B1(_1786_),
    .B2(\third_row[12][3] ),
    .X(_2361_));
 sky130_fd_sc_hd__a221o_1 _4435_ (.A1(\third_row[5][3] ),
    .A2(_1951_),
    .B1(_1939_),
    .B2(\third_row[3][3] ),
    .C1(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__or3_2 _4436_ (.A(_2358_),
    .B(_2360_),
    .C(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__o22a_1 _4437_ (.A1(\third_row[0][3] ),
    .A2(_1904_),
    .B1(_2356_),
    .B2(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__a221o_1 _4438_ (.A1(\second_row[15][3] ),
    .A2(_1726_),
    .B1(_1933_),
    .B2(\second_row[17][3] ),
    .C1(_1866_),
    .X(_2365_));
 sky130_fd_sc_hd__a22o_1 _4439_ (.A1(\second_row[8][3] ),
    .A2(_1828_),
    .B1(_1877_),
    .B2(\second_row[1][3] ),
    .X(_2366_));
 sky130_fd_sc_hd__a221o_1 _4440_ (.A1(\second_row[11][3] ),
    .A2(_1799_),
    .B1(_1868_),
    .B2(\second_row[2][3] ),
    .C1(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__a22o_1 _4441_ (.A1(\second_row[6][3] ),
    .A2(_1831_),
    .B1(_1803_),
    .B2(\second_row[10][3] ),
    .X(_2368_));
 sky130_fd_sc_hd__a221o_1 _4442_ (.A1(\second_row[7][3] ),
    .A2(_1906_),
    .B1(_1911_),
    .B2(\second_row[14][3] ),
    .C1(_2368_),
    .X(_2369_));
 sky130_fd_sc_hd__a22o_1 _4443_ (.A1(\second_row[12][3] ),
    .A2(_1817_),
    .B1(_1785_),
    .B2(\second_row[13][3] ),
    .X(_2370_));
 sky130_fd_sc_hd__a221o_1 _4444_ (.A1(\second_row[16][3] ),
    .A2(_1923_),
    .B1(_1939_),
    .B2(\second_row[4][3] ),
    .C1(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__and3_1 _4445_ (.A(\second_row[9][3] ),
    .B(_1853_),
    .C(_1796_),
    .X(_2372_));
 sky130_fd_sc_hd__a221o_1 _4446_ (.A1(\second_row[3][3] ),
    .A2(_1936_),
    .B1(_1914_),
    .B2(\second_row[5][3] ),
    .C1(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__or4_1 _4447_ (.A(_2367_),
    .B(_2369_),
    .C(_2371_),
    .D(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__o22a_1 _4448_ (.A1(\second_row[0][3] ),
    .A2(_1865_),
    .B1(_2365_),
    .B2(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__xor2_2 _4449_ (.A(_2364_),
    .B(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__nor3_1 _4450_ (.A(_2276_),
    .B(_2286_),
    .C(_2297_),
    .Y(_2377_));
 sky130_fd_sc_hd__and2_1 _4451_ (.A(_2364_),
    .B(_2375_),
    .X(_2378_));
 sky130_fd_sc_hd__a211o_1 _4452_ (.A1(_2353_),
    .A2(_2376_),
    .B1(_2377_),
    .C1(_2378_),
    .X(_2379_));
 sky130_fd_sc_hd__nor3_1 _4453_ (.A(_2253_),
    .B(_2263_),
    .C(_2274_),
    .Y(_2380_));
 sky130_fd_sc_hd__a31o_1 _4454_ (.A1(_2275_),
    .A2(_2298_),
    .A3(_2379_),
    .B1(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__a22o_1 _4455_ (.A1(\third_row[8][6] ),
    .A2(_1955_),
    .B1(_1945_),
    .B2(\third_row[10][6] ),
    .X(_2382_));
 sky130_fd_sc_hd__a221o_1 _4456_ (.A1(\third_row[13][6] ),
    .A2(_1912_),
    .B1(_1949_),
    .B2(\third_row[12][6] ),
    .C1(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__a22o_1 _4457_ (.A1(\third_row[6][6] ),
    .A2(_1907_),
    .B1(_1909_),
    .B2(\third_row[9][6] ),
    .X(_2384_));
 sky130_fd_sc_hd__a221o_1 _4458_ (.A1(\third_row[14][6] ),
    .A2(_1727_),
    .B1(_1915_),
    .B2(\third_row[4][6] ),
    .C1(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__a22o_1 _4459_ (.A1(\third_row[15][6] ),
    .A2(_1923_),
    .B1(_1929_),
    .B2(\third_row[1][6] ),
    .X(_2386_));
 sky130_fd_sc_hd__a221o_1 _4460_ (.A1(\third_row[11][6] ),
    .A2(_1927_),
    .B1(_1921_),
    .B2(\third_row[7][6] ),
    .C1(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__a22o_1 _4461_ (.A1(\third_row[2][6] ),
    .A2(_1937_),
    .B1(_1939_),
    .B2(\third_row[3][6] ),
    .X(_2388_));
 sky130_fd_sc_hd__a221o_1 _4462_ (.A1(\third_row[5][6] ),
    .A2(_1952_),
    .B1(_1943_),
    .B2(\third_row[17][6] ),
    .C1(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__a2111o_1 _4463_ (.A1(\third_row[16][6] ),
    .A2(_1934_),
    .B1(_1919_),
    .C1(_2387_),
    .D1(_2389_),
    .X(_2390_));
 sky130_fd_sc_hd__o32a_2 _4464_ (.A1(_2383_),
    .A2(_2385_),
    .A3(_2390_),
    .B1(_1904_),
    .B2(\third_row[0][6] ),
    .X(_2391_));
 sky130_fd_sc_hd__a221o_1 _4465_ (.A1(\second_row[15][6] ),
    .A2(_1727_),
    .B1(_1934_),
    .B2(\second_row[17][6] ),
    .C1(_1866_),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _4466_ (.A1(\second_row[4][6] ),
    .A2(_1940_),
    .B1(_1877_),
    .B2(\second_row[1][6] ),
    .X(_2393_));
 sky130_fd_sc_hd__a221o_1 _4467_ (.A1(\second_row[5][6] ),
    .A2(_1915_),
    .B1(_1909_),
    .B2(\second_row[10][6] ),
    .C1(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__a22o_1 _4468_ (.A1(\second_row[16][6] ),
    .A2(_1924_),
    .B1(_1929_),
    .B2(\second_row[2][6] ),
    .X(_2395_));
 sky130_fd_sc_hd__a22o_1 _4469_ (.A1(\second_row[3][6] ),
    .A2(_1936_),
    .B1(_1786_),
    .B2(\second_row[13][6] ),
    .X(_2396_));
 sky130_fd_sc_hd__a221o_1 _4470_ (.A1(\second_row[9][6] ),
    .A2(_1955_),
    .B1(_1921_),
    .B2(\second_row[8][6] ),
    .C1(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__a22o_1 _4471_ (.A1(\second_row[6][6] ),
    .A2(_1951_),
    .B1(_1911_),
    .B2(\second_row[14][6] ),
    .X(_2398_));
 sky130_fd_sc_hd__a221o_1 _4472_ (.A1(\second_row[7][6] ),
    .A2(_1906_),
    .B1(_1927_),
    .B2(\second_row[12][6] ),
    .C1(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__a2111o_1 _4473_ (.A1(\second_row[11][6] ),
    .A2(_1946_),
    .B1(_2395_),
    .C1(_2397_),
    .D1(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__o32a_1 _4474_ (.A1(_2392_),
    .A2(_2394_),
    .A3(_2400_),
    .B1(_1865_),
    .B2(\second_row[0][6] ),
    .X(_2401_));
 sky130_fd_sc_hd__or2_1 _4475_ (.A(_2391_),
    .B(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__and2_1 _4476_ (.A(_2391_),
    .B(_2401_),
    .X(_2403_));
 sky130_fd_sc_hd__a21o_1 _4477_ (.A1(_2381_),
    .A2(_2402_),
    .B1(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__nor2_1 _4478_ (.A(_2252_),
    .B(_2404_),
    .Y(_2405_));
 sky130_fd_sc_hd__o22ai_1 _4479_ (.A1(_2068_),
    .A2(_2228_),
    .B1(_2251_),
    .B2(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__nor2_1 _4480_ (.A(_2068_),
    .B(_2069_),
    .Y(_2407_));
 sky130_fd_sc_hd__xnor2_1 _4481_ (.A(_2227_),
    .B(_2407_),
    .Y(_2408_));
 sky130_fd_sc_hd__nor2_1 _4482_ (.A(_2251_),
    .B(_2252_),
    .Y(_2409_));
 sky130_fd_sc_hd__xnor2_1 _4483_ (.A(_2404_),
    .B(_2409_),
    .Y(_2410_));
 sky130_fd_sc_hd__or2_1 _4484_ (.A(_2408_),
    .B(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__and2b_1 _4485_ (.A_N(_2226_),
    .B(_2225_),
    .X(_2412_));
 sky130_fd_sc_hd__xnor2_1 _4486_ (.A(_2202_),
    .B(_2412_),
    .Y(_2413_));
 sky130_fd_sc_hd__and2b_1 _4487_ (.A_N(_2403_),
    .B(_2402_),
    .X(_2414_));
 sky130_fd_sc_hd__xnor2_1 _4488_ (.A(_2381_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__or2_1 _4489_ (.A(_2413_),
    .B(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__and2b_1 _4490_ (.A_N(_2380_),
    .B(_2275_),
    .X(_2417_));
 sky130_fd_sc_hd__nand3_1 _4491_ (.A(_2298_),
    .B(_2379_),
    .C(_2417_),
    .Y(_2418_));
 sky130_fd_sc_hd__or2b_1 _4492_ (.A(_2201_),
    .B_N(_2092_),
    .X(_2419_));
 sky130_fd_sc_hd__xnor2_1 _4493_ (.A(_2200_),
    .B(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__a21o_1 _4494_ (.A1(_2298_),
    .A2(_2379_),
    .B1(_2417_),
    .X(_2421_));
 sky130_fd_sc_hd__nand3_1 _4495_ (.A(_2418_),
    .B(_2420_),
    .C(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__nand2_1 _4496_ (.A(_2140_),
    .B(_2197_),
    .Y(_2423_));
 sky130_fd_sc_hd__xnor2_1 _4497_ (.A(_2115_),
    .B(_2198_),
    .Y(_2424_));
 sky130_fd_sc_hd__xnor2_1 _4498_ (.A(_2423_),
    .B(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__a21oi_1 _4499_ (.A1(_2353_),
    .A2(_2376_),
    .B1(_2378_),
    .Y(_2426_));
 sky130_fd_sc_hd__inv_2 _4500_ (.A(_2298_),
    .Y(_2427_));
 sky130_fd_sc_hd__nor2_1 _4501_ (.A(_2427_),
    .B(_2377_),
    .Y(_2428_));
 sky130_fd_sc_hd__xnor2_1 _4502_ (.A(_2426_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__nand2_1 _4503_ (.A(_2425_),
    .B(_2429_),
    .Y(_2430_));
 sky130_fd_sc_hd__xnor2_1 _4504_ (.A(_2353_),
    .B(_2376_),
    .Y(_2431_));
 sky130_fd_sc_hd__a21o_1 _4505_ (.A1(_2171_),
    .A2(_2194_),
    .B1(_2196_),
    .X(_2432_));
 sky130_fd_sc_hd__or4_1 _4506_ (.A(_2117_),
    .B(_2128_),
    .C(_2129_),
    .D(_2139_),
    .X(_2433_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_2140_),
    .B(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__xnor2_1 _4508_ (.A(_2432_),
    .B(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__and2b_1 _4509_ (.A_N(_2431_),
    .B(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__inv_2 _4510_ (.A(_2436_),
    .Y(_2437_));
 sky130_fd_sc_hd__xor2_1 _4511_ (.A(_2431_),
    .B(_2435_),
    .X(_2438_));
 sky130_fd_sc_hd__xor2_1 _4512_ (.A(_2328_),
    .B(_2351_),
    .X(_2439_));
 sky130_fd_sc_hd__xor2_1 _4513_ (.A(_2171_),
    .B(_2194_),
    .X(_2440_));
 sky130_fd_sc_hd__xor2_1 _4514_ (.A(_2439_),
    .B(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__xor2_2 _4515_ (.A(_1859_),
    .B(_2170_),
    .X(_2442_));
 sky130_fd_sc_hd__xor2_2 _4516_ (.A(_1897_),
    .B(_2327_),
    .X(_2443_));
 sky130_fd_sc_hd__xor2_2 _4517_ (.A(_2442_),
    .B(_2443_),
    .X(_2444_));
 sky130_fd_sc_hd__a32o_1 _4518_ (.A1(_1862_),
    .A2(_1900_),
    .A3(_2444_),
    .B1(_2443_),
    .B2(_2442_),
    .X(_2445_));
 sky130_fd_sc_hd__and2_1 _4519_ (.A(_2439_),
    .B(_2440_),
    .X(_2446_));
 sky130_fd_sc_hd__a21oi_2 _4520_ (.A1(_2441_),
    .A2(_2445_),
    .B1(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__or2_1 _4521_ (.A(_2438_),
    .B(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__nor2_1 _4522_ (.A(_2425_),
    .B(_2429_),
    .Y(_2449_));
 sky130_fd_sc_hd__a21oi_1 _4523_ (.A1(_2418_),
    .A2(_2421_),
    .B1(_2420_),
    .Y(_2450_));
 sky130_fd_sc_hd__a311o_1 _4524_ (.A1(_2430_),
    .A2(_2437_),
    .A3(_2448_),
    .B1(_2449_),
    .C1(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__and2_1 _4525_ (.A(_2413_),
    .B(_2415_),
    .X(_2452_));
 sky130_fd_sc_hd__a31o_1 _4526_ (.A1(_2416_),
    .A2(_2422_),
    .A3(_2451_),
    .B1(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__and2_1 _4527_ (.A(_2408_),
    .B(_2410_),
    .X(_2454_));
 sky130_fd_sc_hd__a21oi_1 _4528_ (.A1(_2411_),
    .A2(_2453_),
    .B1(_2454_),
    .Y(_2455_));
 sky130_fd_sc_hd__nor4_1 _4529_ (.A(_2068_),
    .B(_2228_),
    .C(_2251_),
    .D(_2405_),
    .Y(_2456_));
 sky130_fd_sc_hd__a21o_1 _4530_ (.A1(_2406_),
    .A2(_2455_),
    .B1(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__nor2_1 _4531_ (.A(_2044_),
    .B(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__xor2_1 _4532_ (.A(_2408_),
    .B(_2410_),
    .X(_2459_));
 sky130_fd_sc_hd__xnor2_1 _4533_ (.A(_2453_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_2008_),
    .B(_2019_),
    .Y(_2461_));
 sky130_fd_sc_hd__xnor2_1 _4535_ (.A(_2461_),
    .B(_2030_),
    .Y(_2462_));
 sky130_fd_sc_hd__nor2_1 _4536_ (.A(_2460_),
    .B(_2462_),
    .Y(_2463_));
 sky130_fd_sc_hd__inv_2 _4537_ (.A(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__and2b_1 _4538_ (.A_N(_2007_),
    .B(_1971_),
    .X(_2465_));
 sky130_fd_sc_hd__or2_1 _4539_ (.A(_2008_),
    .B(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__o21ba_1 _4540_ (.A1(_2438_),
    .A2(_2447_),
    .B1_N(_2436_),
    .X(_2467_));
 sky130_fd_sc_hd__o21a_1 _4541_ (.A1(_2449_),
    .A2(_2467_),
    .B1(_2430_),
    .X(_2468_));
 sky130_fd_sc_hd__and3_1 _4542_ (.A(_2418_),
    .B(_2420_),
    .C(_2421_),
    .X(_2469_));
 sky130_fd_sc_hd__nor2_1 _4543_ (.A(_2469_),
    .B(_2450_),
    .Y(_2470_));
 sky130_fd_sc_hd__xor2_1 _4544_ (.A(_2468_),
    .B(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__xor2_1 _4545_ (.A(_2466_),
    .B(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__xnor2_1 _4546_ (.A(_2438_),
    .B(_2447_),
    .Y(_2473_));
 sky130_fd_sc_hd__nor3_1 _4547_ (.A(_2005_),
    .B(_1983_),
    .C(_1994_),
    .Y(_2474_));
 sky130_fd_sc_hd__nor2_1 _4548_ (.A(_2006_),
    .B(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__xnor2_1 _4549_ (.A(_2473_),
    .B(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__xor2_1 _4550_ (.A(_2441_),
    .B(_2445_),
    .X(_2477_));
 sky130_fd_sc_hd__and2b_1 _4551_ (.A_N(_2005_),
    .B(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__and2b_1 _4552_ (.A_N(_2473_),
    .B(_2475_),
    .X(_2479_));
 sky130_fd_sc_hd__a21o_1 _4553_ (.A1(_2476_),
    .A2(_2478_),
    .B1(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__and2b_1 _4554_ (.A_N(_2006_),
    .B(_1982_),
    .X(_2481_));
 sky130_fd_sc_hd__or2_1 _4555_ (.A(_2007_),
    .B(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__xnor2_1 _4556_ (.A(_2425_),
    .B(_2429_),
    .Y(_2483_));
 sky130_fd_sc_hd__xnor2_1 _4557_ (.A(_2467_),
    .B(_2483_),
    .Y(_2484_));
 sky130_fd_sc_hd__xor2_1 _4558_ (.A(_2482_),
    .B(_2484_),
    .X(_2485_));
 sky130_fd_sc_hd__nor2_1 _4559_ (.A(_2482_),
    .B(_2484_),
    .Y(_2486_));
 sky130_fd_sc_hd__a21o_1 _4560_ (.A1(_2480_),
    .A2(_2485_),
    .B1(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__nor2_1 _4561_ (.A(_2466_),
    .B(_2471_),
    .Y(_2488_));
 sky130_fd_sc_hd__a21o_1 _4562_ (.A1(_2472_),
    .A2(_2487_),
    .B1(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__xnor2_2 _4563_ (.A(_2008_),
    .B(_2019_),
    .Y(_2490_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_2422_),
    .B(_2451_),
    .Y(_2491_));
 sky130_fd_sc_hd__or2b_1 _4565_ (.A(_2452_),
    .B_N(_2416_),
    .X(_2492_));
 sky130_fd_sc_hd__xor2_2 _4566_ (.A(_2491_),
    .B(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__xor2_2 _4567_ (.A(_2490_),
    .B(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__and2_1 _4568_ (.A(_2460_),
    .B(_2462_),
    .X(_2495_));
 sky130_fd_sc_hd__nor2_1 _4569_ (.A(_2490_),
    .B(_2493_),
    .Y(_2496_));
 sky130_fd_sc_hd__a211o_1 _4570_ (.A1(_2489_),
    .A2(_2494_),
    .B1(_2495_),
    .C1(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__xor2_1 _4571_ (.A(_2031_),
    .B(_1960_),
    .X(_2498_));
 sky130_fd_sc_hd__and2b_1 _4572_ (.A_N(_2456_),
    .B(_2406_),
    .X(_2499_));
 sky130_fd_sc_hd__xnor2_1 _4573_ (.A(_2455_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_2498_),
    .B(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hd__and2_1 _4575_ (.A(_2044_),
    .B(_2457_),
    .X(_2502_));
 sky130_fd_sc_hd__nor2_1 _4576_ (.A(_2498_),
    .B(_2500_),
    .Y(_2503_));
 sky130_fd_sc_hd__a311oi_1 _4577_ (.A1(_2464_),
    .A2(_2497_),
    .A3(_2501_),
    .B1(_2502_),
    .C1(_2503_),
    .Y(_2504_));
 sky130_fd_sc_hd__or3b_1 _4578_ (.A(_1960_),
    .B(_2043_),
    .C_N(_2031_),
    .X(_2505_));
 sky130_fd_sc_hd__o21a_2 _4579_ (.A1(_2458_),
    .A2(_2504_),
    .B1(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__xor2_1 _4580_ (.A(_1901_),
    .B(_2444_),
    .X(_2507_));
 sky130_fd_sc_hd__or2_1 _4581_ (.A(_1903_),
    .B(_2507_),
    .X(_2508_));
 sky130_fd_sc_hd__xor2_1 _4582_ (.A(_2005_),
    .B(_2477_),
    .X(_2509_));
 sky130_fd_sc_hd__or2b_1 _4583_ (.A(_2508_),
    .B_N(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__xnor2_1 _4584_ (.A(_2476_),
    .B(_2478_),
    .Y(_2511_));
 sky130_fd_sc_hd__or2b_1 _4585_ (.A(_2510_),
    .B_N(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__xnor2_1 _4586_ (.A(_2480_),
    .B(_2485_),
    .Y(_2513_));
 sky130_fd_sc_hd__or2b_1 _4587_ (.A(_2512_),
    .B_N(_2513_),
    .X(_2514_));
 sky130_fd_sc_hd__xnor2_1 _4588_ (.A(_2472_),
    .B(_2487_),
    .Y(_2515_));
 sky130_fd_sc_hd__or2b_1 _4589_ (.A(_2514_),
    .B_N(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__xnor2_2 _4590_ (.A(_2489_),
    .B(_2494_),
    .Y(_2517_));
 sky130_fd_sc_hd__or2b_1 _4591_ (.A(_2516_),
    .B_N(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__a21o_1 _4592_ (.A1(_2489_),
    .A2(_2494_),
    .B1(_2496_),
    .X(_2519_));
 sky130_fd_sc_hd__nor2_1 _4593_ (.A(_2463_),
    .B(_2495_),
    .Y(_2520_));
 sky130_fd_sc_hd__xnor2_1 _4594_ (.A(_2519_),
    .B(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__or2b_1 _4595_ (.A(_2518_),
    .B_N(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__nor2_1 _4596_ (.A(_2458_),
    .B(_2502_),
    .Y(_2523_));
 sky130_fd_sc_hd__a31o_1 _4597_ (.A1(_2464_),
    .A2(_2497_),
    .A3(_2501_),
    .B1(_2503_),
    .X(_2524_));
 sky130_fd_sc_hd__xnor2_2 _4598_ (.A(_2523_),
    .B(_2524_),
    .Y(_2525_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_2464_),
    .B(_2497_),
    .Y(_2526_));
 sky130_fd_sc_hd__and2b_1 _4600_ (.A_N(_2503_),
    .B(_2501_),
    .X(_2527_));
 sky130_fd_sc_hd__xor2_2 _4601_ (.A(_2526_),
    .B(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__a22oi_4 _4602_ (.A1(_2506_),
    .A2(_2522_),
    .B1(_2525_),
    .B2(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__o211a_2 _4603_ (.A1(_2525_),
    .A2(_2528_),
    .B1(_2506_),
    .C1(_2522_),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_8 _4604_ (.A(net9),
    .X(_2531_));
 sky130_fd_sc_hd__inv_2 _4605_ (.A(_2531_),
    .Y(_0000_));
 sky130_fd_sc_hd__o31a_1 _4606_ (.A1(_1903_),
    .A2(_2529_),
    .A3(_2530_),
    .B1(_0000_),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 _4607_ (.A(_2506_),
    .X(_2532_));
 sky130_fd_sc_hd__a21boi_1 _4608_ (.A1(_1903_),
    .A2(_2532_),
    .B1_N(_2507_),
    .Y(_2533_));
 sky130_fd_sc_hd__and3b_1 _4609_ (.A_N(_2444_),
    .B(_2506_),
    .C(_1903_),
    .X(_2534_));
 sky130_fd_sc_hd__o41a_1 _4610_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2533_),
    .A4(_2534_),
    .B1(_0000_),
    .X(net12));
 sky130_fd_sc_hd__a21oi_1 _4611_ (.A1(_2532_),
    .A2(_2508_),
    .B1(_2509_),
    .Y(_2535_));
 sky130_fd_sc_hd__and3_1 _4612_ (.A(_2532_),
    .B(_2509_),
    .C(_2508_),
    .X(_2536_));
 sky130_fd_sc_hd__o41a_1 _4613_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2535_),
    .A4(_2536_),
    .B1(_0000_),
    .X(net13));
 sky130_fd_sc_hd__a21oi_1 _4614_ (.A1(_2532_),
    .A2(_2510_),
    .B1(_2511_),
    .Y(_2537_));
 sky130_fd_sc_hd__and3_1 _4615_ (.A(_2532_),
    .B(_2511_),
    .C(_2510_),
    .X(_2538_));
 sky130_fd_sc_hd__o41a_1 _4616_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2537_),
    .A4(_2538_),
    .B1(_0000_),
    .X(net14));
 sky130_fd_sc_hd__a21oi_1 _4617_ (.A1(_2532_),
    .A2(_2512_),
    .B1(_2513_),
    .Y(_2539_));
 sky130_fd_sc_hd__and3_1 _4618_ (.A(_2532_),
    .B(_2513_),
    .C(_2512_),
    .X(_2540_));
 sky130_fd_sc_hd__o41a_1 _4619_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2539_),
    .A4(_2540_),
    .B1(_0000_),
    .X(net15));
 sky130_fd_sc_hd__a21oi_1 _4620_ (.A1(_2532_),
    .A2(_2514_),
    .B1(_2515_),
    .Y(_2541_));
 sky130_fd_sc_hd__and3_1 _4621_ (.A(_2506_),
    .B(_2514_),
    .C(_2515_),
    .X(_2542_));
 sky130_fd_sc_hd__o41a_1 _4622_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2541_),
    .A4(_2542_),
    .B1(_0000_),
    .X(net16));
 sky130_fd_sc_hd__a21oi_1 _4623_ (.A1(_2532_),
    .A2(_2516_),
    .B1(_2517_),
    .Y(_2543_));
 sky130_fd_sc_hd__and3_1 _4624_ (.A(_2506_),
    .B(_2516_),
    .C(_2517_),
    .X(_2544_));
 sky130_fd_sc_hd__o41a_1 _4625_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2543_),
    .A4(_2544_),
    .B1(_0000_),
    .X(net17));
 sky130_fd_sc_hd__a21oi_1 _4626_ (.A1(_2532_),
    .A2(_2518_),
    .B1(_2521_),
    .Y(_2545_));
 sky130_fd_sc_hd__and3_1 _4627_ (.A(_2506_),
    .B(_2518_),
    .C(_2521_),
    .X(_2546_));
 sky130_fd_sc_hd__o41a_1 _4628_ (.A1(_2529_),
    .A2(_2530_),
    .A3(_2545_),
    .A4(_2546_),
    .B1(_0000_),
    .X(net18));
 sky130_fd_sc_hd__a21oi_1 _4629_ (.A1(_1067_),
    .A2(_1607_),
    .B1(net9),
    .Y(_2547_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(net19),
    .A1(_1617_),
    .S(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_1 _4631_ (.A(_2548_),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_8 _4632_ (.A(_2531_),
    .X(_2549_));
 sky130_fd_sc_hd__buf_4 _4633_ (.A(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__inv_2 _4634_ (.A(_2550_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _4635_ (.A(_2550_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(_2550_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _4637_ (.A(_2550_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _4638_ (.A(_2550_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _4639_ (.A(_2550_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _4640_ (.A(_2550_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _4641_ (.A(_2550_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _4642_ (.A(_2550_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _4643_ (.A(_2550_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_4 _4644_ (.A(_2549_),
    .X(_2551_));
 sky130_fd_sc_hd__inv_2 _4645_ (.A(_2551_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _4646_ (.A(_2551_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _4647_ (.A(_2551_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(_2551_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _4649_ (.A(_2551_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _4650_ (.A(_2551_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _4651_ (.A(_2551_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _4652_ (.A(_2551_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _4653_ (.A(_2551_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _4654_ (.A(_2551_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_4 _4655_ (.A(_2549_),
    .X(_2552_));
 sky130_fd_sc_hd__inv_2 _4656_ (.A(_2552_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _4657_ (.A(_2552_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _4658_ (.A(_2552_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _4659_ (.A(_2552_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _4660_ (.A(_2552_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _4661_ (.A(_2552_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _4662_ (.A(_2552_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _4663_ (.A(_2552_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _4664_ (.A(_2552_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _4665_ (.A(_2552_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_4 _4666_ (.A(_2549_),
    .X(_2553_));
 sky130_fd_sc_hd__inv_2 _4667_ (.A(_2553_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _4668_ (.A(_2553_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _4669_ (.A(_2553_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _4670_ (.A(_2553_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _4671_ (.A(_2553_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _4672_ (.A(_2553_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _4673_ (.A(_2553_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _4674_ (.A(_2553_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _4675_ (.A(_2553_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _4676_ (.A(_2553_),
    .Y(_0040_));
 sky130_fd_sc_hd__buf_4 _4677_ (.A(_2549_),
    .X(_2554_));
 sky130_fd_sc_hd__inv_2 _4678_ (.A(_2554_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _4679_ (.A(_2554_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _4680_ (.A(_2554_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _4681_ (.A(_2554_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _4682_ (.A(_2554_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _4683_ (.A(_2554_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _4684_ (.A(_2554_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _4685_ (.A(_2554_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _4686_ (.A(_2554_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _4687_ (.A(_2554_),
    .Y(_0050_));
 sky130_fd_sc_hd__buf_4 _4688_ (.A(_2549_),
    .X(_2555_));
 sky130_fd_sc_hd__inv_2 _4689_ (.A(_2555_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(_2555_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _4691_ (.A(_2555_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _4692_ (.A(_2555_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _4693_ (.A(_2555_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _4694_ (.A(_2555_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _4695_ (.A(_2555_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _4696_ (.A(_2555_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _4697_ (.A(_2555_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _4698_ (.A(_2555_),
    .Y(_0060_));
 sky130_fd_sc_hd__buf_4 _4699_ (.A(_2549_),
    .X(_2556_));
 sky130_fd_sc_hd__inv_2 _4700_ (.A(_2556_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _4701_ (.A(_2556_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _4702_ (.A(_2556_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _4703_ (.A(_2556_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _4704_ (.A(_2556_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _4705_ (.A(_2556_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _4706_ (.A(_2556_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _4707_ (.A(_2556_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _4708_ (.A(_2556_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _4709_ (.A(_2556_),
    .Y(_0070_));
 sky130_fd_sc_hd__buf_4 _4710_ (.A(_2549_),
    .X(_2557_));
 sky130_fd_sc_hd__inv_2 _4711_ (.A(_2557_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _4712_ (.A(_2557_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _4713_ (.A(_2557_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _4714_ (.A(_2557_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _4715_ (.A(_2557_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _4716_ (.A(_2557_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _4717_ (.A(_2557_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _4718_ (.A(_2557_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _4719_ (.A(_2557_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _4720_ (.A(_2557_),
    .Y(_0080_));
 sky130_fd_sc_hd__buf_4 _4721_ (.A(_2531_),
    .X(_2558_));
 sky130_fd_sc_hd__buf_4 _4722_ (.A(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__inv_2 _4723_ (.A(_2559_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _4724_ (.A(_2559_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _4725_ (.A(_2559_),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _4726_ (.A(_2559_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _4727_ (.A(_2559_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _4728_ (.A(_2559_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _4729_ (.A(_2559_),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _4730_ (.A(_2559_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _4731_ (.A(_2559_),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _4732_ (.A(_2559_),
    .Y(_0090_));
 sky130_fd_sc_hd__buf_4 _4733_ (.A(_2558_),
    .X(_2560_));
 sky130_fd_sc_hd__inv_2 _4734_ (.A(_2560_),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _4735_ (.A(_2560_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _4736_ (.A(_2560_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _4737_ (.A(_2560_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _4738_ (.A(_2560_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _4739_ (.A(_2560_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _4740_ (.A(_2560_),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _4741_ (.A(_2560_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _4742_ (.A(_2560_),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _4743_ (.A(_2560_),
    .Y(_0100_));
 sky130_fd_sc_hd__buf_4 _4744_ (.A(_2558_),
    .X(_2561_));
 sky130_fd_sc_hd__inv_2 _4745_ (.A(_2561_),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _4746_ (.A(_2561_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _4747_ (.A(_2561_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _4748_ (.A(_2561_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _4749_ (.A(_2561_),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _4750_ (.A(_2561_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _4751_ (.A(_2561_),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _4752_ (.A(_2561_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _4753_ (.A(_2561_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _4754_ (.A(_2561_),
    .Y(_0110_));
 sky130_fd_sc_hd__buf_4 _4755_ (.A(_2558_),
    .X(_2562_));
 sky130_fd_sc_hd__inv_2 _4756_ (.A(_2562_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _4757_ (.A(_2562_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _4758_ (.A(_2562_),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _4759_ (.A(_2562_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _4760_ (.A(_2562_),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _4761_ (.A(_2562_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _4762_ (.A(_2562_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _4763_ (.A(_2562_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _4764_ (.A(_2562_),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _4765_ (.A(_2562_),
    .Y(_0120_));
 sky130_fd_sc_hd__clkbuf_8 _4766_ (.A(_2558_),
    .X(_2563_));
 sky130_fd_sc_hd__inv_2 _4767_ (.A(_2563_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _4768_ (.A(_2563_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _4769_ (.A(_2563_),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _4770_ (.A(_2563_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _4771_ (.A(_2563_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _4772_ (.A(_2563_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _4773_ (.A(_2563_),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _4774_ (.A(_2563_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _4775_ (.A(_2563_),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _4776_ (.A(_2563_),
    .Y(_0130_));
 sky130_fd_sc_hd__buf_4 _4777_ (.A(_2558_),
    .X(_2564_));
 sky130_fd_sc_hd__inv_2 _4778_ (.A(_2564_),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _4779_ (.A(_2564_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _4780_ (.A(_2564_),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _4781_ (.A(_2564_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _4782_ (.A(_2564_),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _4783_ (.A(_2564_),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _4784_ (.A(_2564_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _4785_ (.A(_2564_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _4786_ (.A(_2564_),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _4787_ (.A(_2564_),
    .Y(_0140_));
 sky130_fd_sc_hd__clkbuf_8 _4788_ (.A(_2558_),
    .X(_2565_));
 sky130_fd_sc_hd__inv_2 _4789_ (.A(_2565_),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _4790_ (.A(_2565_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _4791_ (.A(_2565_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _4792_ (.A(_2565_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _4793_ (.A(_2565_),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _4794_ (.A(_2565_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _4795_ (.A(_2565_),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _4796_ (.A(_2565_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _4797_ (.A(_2565_),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _4798_ (.A(_2565_),
    .Y(_0150_));
 sky130_fd_sc_hd__buf_4 _4799_ (.A(_2558_),
    .X(_2566_));
 sky130_fd_sc_hd__inv_2 _4800_ (.A(_2566_),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _4801_ (.A(_2566_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _4802_ (.A(_2566_),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _4803_ (.A(_2566_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _4804_ (.A(_2566_),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _4805_ (.A(_2566_),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _4806_ (.A(_2566_),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _4807_ (.A(_2566_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _4808_ (.A(_2566_),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _4809_ (.A(_2566_),
    .Y(_0160_));
 sky130_fd_sc_hd__clkbuf_8 _4810_ (.A(_2558_),
    .X(_2567_));
 sky130_fd_sc_hd__inv_2 _4811_ (.A(_2567_),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _4812_ (.A(_2567_),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _4813_ (.A(_2567_),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _4814_ (.A(_2567_),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _4815_ (.A(_2567_),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _4816_ (.A(_2567_),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _4817_ (.A(_2567_),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _4818_ (.A(_2567_),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _4819_ (.A(_2567_),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _4820_ (.A(_2567_),
    .Y(_0170_));
 sky130_fd_sc_hd__clkbuf_8 _4821_ (.A(_2558_),
    .X(_2568_));
 sky130_fd_sc_hd__inv_2 _4822_ (.A(_2568_),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _4823_ (.A(_2568_),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _4824_ (.A(_2568_),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4825_ (.A(_2568_),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _4826_ (.A(_2568_),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _4827_ (.A(_2568_),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _4828_ (.A(_2568_),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _4829_ (.A(_2568_),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _4830_ (.A(_2568_),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _4831_ (.A(_2568_),
    .Y(_0180_));
 sky130_fd_sc_hd__clkbuf_4 _4832_ (.A(_2531_),
    .X(_2569_));
 sky130_fd_sc_hd__buf_4 _4833_ (.A(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__inv_2 _4834_ (.A(_2570_),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _4835_ (.A(_2570_),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _4836_ (.A(_2570_),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _4837_ (.A(_2570_),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _4838_ (.A(_2570_),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _4839_ (.A(_2570_),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _4840_ (.A(_2570_),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _4841_ (.A(_2570_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _4842_ (.A(_2570_),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _4843_ (.A(_2570_),
    .Y(_0190_));
 sky130_fd_sc_hd__clkbuf_8 _4844_ (.A(_2569_),
    .X(_2571_));
 sky130_fd_sc_hd__inv_2 _4845_ (.A(_2571_),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _4846_ (.A(_2571_),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _4847_ (.A(_2571_),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _4848_ (.A(_2571_),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _4849_ (.A(_2571_),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _4850_ (.A(_2571_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _4851_ (.A(_2571_),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _4852_ (.A(_2571_),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _4853_ (.A(_2571_),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _4854_ (.A(_2571_),
    .Y(_0200_));
 sky130_fd_sc_hd__buf_4 _4855_ (.A(_2569_),
    .X(_2572_));
 sky130_fd_sc_hd__inv_2 _4856_ (.A(_2572_),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _4857_ (.A(_2572_),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _4858_ (.A(_2572_),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _4859_ (.A(_2572_),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _4860_ (.A(_2572_),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _4861_ (.A(_2572_),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _4862_ (.A(_2572_),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _4863_ (.A(_2572_),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _4864_ (.A(_2572_),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _4865_ (.A(_2572_),
    .Y(_0210_));
 sky130_fd_sc_hd__buf_4 _4866_ (.A(_2569_),
    .X(_2573_));
 sky130_fd_sc_hd__inv_2 _4867_ (.A(_2573_),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _4868_ (.A(_2573_),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _4869_ (.A(_2573_),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _4870_ (.A(_2573_),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _4871_ (.A(_2573_),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _4872_ (.A(_2573_),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _4873_ (.A(_2573_),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _4874_ (.A(_2573_),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _4875_ (.A(_2573_),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _4876_ (.A(_2573_),
    .Y(_0220_));
 sky130_fd_sc_hd__buf_4 _4877_ (.A(_2569_),
    .X(_2574_));
 sky130_fd_sc_hd__inv_2 _4878_ (.A(_2574_),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _4879_ (.A(_2574_),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _4880_ (.A(_2574_),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _4881_ (.A(_2574_),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _4882_ (.A(_2574_),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _4883_ (.A(_2574_),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _4884_ (.A(_2574_),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _4885_ (.A(_2574_),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _4886_ (.A(_2574_),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _4887_ (.A(_2574_),
    .Y(_0230_));
 sky130_fd_sc_hd__clkbuf_8 _4888_ (.A(_2569_),
    .X(_2575_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(_2575_),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _4890_ (.A(_2575_),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _4891_ (.A(_2575_),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _4892_ (.A(_2575_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _4893_ (.A(_2575_),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _4894_ (.A(_2575_),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _4895_ (.A(_2575_),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _4896_ (.A(_2575_),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _4897_ (.A(_2575_),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _4898_ (.A(_2575_),
    .Y(_0240_));
 sky130_fd_sc_hd__clkbuf_8 _4899_ (.A(_2569_),
    .X(_2576_));
 sky130_fd_sc_hd__inv_2 _4900_ (.A(_2576_),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _4901_ (.A(_2576_),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _4902_ (.A(_2576_),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _4903_ (.A(_2576_),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _4904_ (.A(_2576_),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _4905_ (.A(_2576_),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _4906_ (.A(_2576_),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _4907_ (.A(_2576_),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _4908_ (.A(_2576_),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _4909_ (.A(_2576_),
    .Y(_0250_));
 sky130_fd_sc_hd__buf_4 _4910_ (.A(_2569_),
    .X(_2577_));
 sky130_fd_sc_hd__inv_2 _4911_ (.A(_2577_),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _4912_ (.A(_2577_),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _4913_ (.A(_2577_),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _4914_ (.A(_2577_),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _4915_ (.A(_2577_),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _4916_ (.A(_2577_),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _4917_ (.A(_2577_),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _4918_ (.A(_2577_),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _4919_ (.A(_2577_),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _4920_ (.A(_2577_),
    .Y(_0260_));
 sky130_fd_sc_hd__clkbuf_8 _4921_ (.A(_2569_),
    .X(_2578_));
 sky130_fd_sc_hd__inv_2 _4922_ (.A(_2578_),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _4923_ (.A(_2578_),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _4924_ (.A(_2578_),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _4925_ (.A(_2578_),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _4926_ (.A(_2578_),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_2 _4927_ (.A(_2578_),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _4928_ (.A(_2578_),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(_2578_),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_2 _4930_ (.A(_2578_),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _4931_ (.A(_2578_),
    .Y(_0270_));
 sky130_fd_sc_hd__clkbuf_8 _4932_ (.A(_2569_),
    .X(_2579_));
 sky130_fd_sc_hd__inv_2 _4933_ (.A(_2579_),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _4934_ (.A(_2579_),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_2 _4935_ (.A(_2579_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _4936_ (.A(_2579_),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_2 _4937_ (.A(_2579_),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _4938_ (.A(_2579_),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _4939_ (.A(_2579_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _4940_ (.A(_2579_),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_2 _4941_ (.A(_2579_),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_2 _4942_ (.A(_2579_),
    .Y(_0280_));
 sky130_fd_sc_hd__buf_4 _4943_ (.A(_2531_),
    .X(_2580_));
 sky130_fd_sc_hd__buf_4 _4944_ (.A(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__inv_2 _4945_ (.A(_2581_),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _4946_ (.A(_2581_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _4947_ (.A(_2581_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _4948_ (.A(_2581_),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_2 _4949_ (.A(_2581_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _4950_ (.A(_2581_),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_2 _4951_ (.A(_2581_),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _4952_ (.A(_2581_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _4953_ (.A(_2581_),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_2 _4954_ (.A(_2581_),
    .Y(_0290_));
 sky130_fd_sc_hd__buf_6 _4955_ (.A(_2580_),
    .X(_2582_));
 sky130_fd_sc_hd__inv_2 _4956_ (.A(_2582_),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_2 _4957_ (.A(_2582_),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _4958_ (.A(_2582_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _4959_ (.A(_2582_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _4960_ (.A(_2582_),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _4961_ (.A(_2582_),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_2 _4962_ (.A(_2582_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _4963_ (.A(_2582_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _4964_ (.A(_2582_),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_2 _4965_ (.A(_2582_),
    .Y(_0300_));
 sky130_fd_sc_hd__clkbuf_8 _4966_ (.A(_2580_),
    .X(_2583_));
 sky130_fd_sc_hd__inv_2 _4967_ (.A(_2583_),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _4968_ (.A(_2583_),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_2 _4969_ (.A(_2583_),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _4970_ (.A(_2583_),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _4971_ (.A(_2583_),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _4972_ (.A(_2583_),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _4973_ (.A(_2583_),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _4974_ (.A(_2583_),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_2 _4975_ (.A(_2583_),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _4976_ (.A(_2583_),
    .Y(_0310_));
 sky130_fd_sc_hd__clkbuf_8 _4977_ (.A(_2580_),
    .X(_2584_));
 sky130_fd_sc_hd__inv_2 _4978_ (.A(_2584_),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _4979_ (.A(_2584_),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_2 _4980_ (.A(_2584_),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _4981_ (.A(_2584_),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_2 _4982_ (.A(_2584_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _4983_ (.A(_2584_),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _4984_ (.A(_2584_),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _4985_ (.A(_2584_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _4986_ (.A(_2584_),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_2 _4987_ (.A(_2584_),
    .Y(_0320_));
 sky130_fd_sc_hd__clkbuf_8 _4988_ (.A(_2580_),
    .X(_2585_));
 sky130_fd_sc_hd__inv_2 _4989_ (.A(_2585_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _4990_ (.A(_2585_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _4991_ (.A(_2585_),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _4992_ (.A(_2585_),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _4993_ (.A(_2585_),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _4994_ (.A(_2585_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _4995_ (.A(_2585_),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_2 _4996_ (.A(_2585_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _4997_ (.A(_2585_),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _4998_ (.A(_2585_),
    .Y(_0330_));
 sky130_fd_sc_hd__clkbuf_8 _4999_ (.A(_2580_),
    .X(_2586_));
 sky130_fd_sc_hd__inv_2 _5000_ (.A(_2586_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _5001_ (.A(_2586_),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _5002_ (.A(_2586_),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _5003_ (.A(_2586_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _5004_ (.A(_2586_),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _5005_ (.A(_2586_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _5006_ (.A(_2586_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _5007_ (.A(_2586_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _5008_ (.A(_2586_),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_2 _5009_ (.A(_2586_),
    .Y(_0340_));
 sky130_fd_sc_hd__clkbuf_8 _5010_ (.A(_2580_),
    .X(_2587_));
 sky130_fd_sc_hd__inv_2 _5011_ (.A(_2587_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _5012_ (.A(_2587_),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_2 _5013_ (.A(_2587_),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_2 _5014_ (.A(_2587_),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _5015_ (.A(_2587_),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _5016_ (.A(_2587_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _5017_ (.A(_2587_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _5018_ (.A(_2587_),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _5019_ (.A(_2587_),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _5020_ (.A(_2587_),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_8 _5021_ (.A(_2580_),
    .X(_2588_));
 sky130_fd_sc_hd__inv_2 _5022_ (.A(_2588_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _5023_ (.A(_2588_),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _5024_ (.A(_2588_),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _5025_ (.A(_2588_),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _5026_ (.A(_2588_),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _5027_ (.A(_2588_),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _5028_ (.A(_2588_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _5029_ (.A(_2588_),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_2 _5030_ (.A(_2588_),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_2 _5031_ (.A(_2588_),
    .Y(_0360_));
 sky130_fd_sc_hd__buf_4 _5032_ (.A(_2580_),
    .X(_2589_));
 sky130_fd_sc_hd__inv_2 _5033_ (.A(_2589_),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _5034_ (.A(_2589_),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _5035_ (.A(_2589_),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_2 _5036_ (.A(_2589_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _5037_ (.A(_2589_),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _5038_ (.A(_2589_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _5039_ (.A(_2589_),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_2 _5040_ (.A(_2589_),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _5041_ (.A(_2589_),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_2 _5042_ (.A(_2589_),
    .Y(_0370_));
 sky130_fd_sc_hd__buf_4 _5043_ (.A(_2580_),
    .X(_2590_));
 sky130_fd_sc_hd__inv_2 _5044_ (.A(_2590_),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_2 _5045_ (.A(_2590_),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _5046_ (.A(_2590_),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_2 _5047_ (.A(_2590_),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_2 _5048_ (.A(_2590_),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_2 _5049_ (.A(_2590_),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _5050_ (.A(_2590_),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_2 _5051_ (.A(_2590_),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_2 _5052_ (.A(_2590_),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_2 _5053_ (.A(_2590_),
    .Y(_0380_));
 sky130_fd_sc_hd__clkbuf_4 _5054_ (.A(net9),
    .X(_2591_));
 sky130_fd_sc_hd__buf_8 _5055_ (.A(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__inv_2 _5056_ (.A(_2592_),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _5057_ (.A(_2592_),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_2 _5058_ (.A(_2592_),
    .Y(_0383_));
 sky130_fd_sc_hd__inv_2 _5059_ (.A(_2592_),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _5060_ (.A(_2592_),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_2 _5061_ (.A(_2592_),
    .Y(_0386_));
 sky130_fd_sc_hd__inv_2 _5062_ (.A(_2592_),
    .Y(_0387_));
 sky130_fd_sc_hd__inv_2 _5063_ (.A(_2592_),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_2 _5064_ (.A(_2592_),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _5065_ (.A(_2592_),
    .Y(_0390_));
 sky130_fd_sc_hd__clkbuf_8 _5066_ (.A(_2591_),
    .X(_2593_));
 sky130_fd_sc_hd__inv_2 _5067_ (.A(_2593_),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _5068_ (.A(_2593_),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_2 _5069_ (.A(_2593_),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_2 _5070_ (.A(_2593_),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_2 _5071_ (.A(_2593_),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_2 _5072_ (.A(_2593_),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_2 _5073_ (.A(_2593_),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_2 _5074_ (.A(_2593_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _5075_ (.A(_2593_),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_2 _5076_ (.A(_2593_),
    .Y(_0400_));
 sky130_fd_sc_hd__clkbuf_8 _5077_ (.A(_2591_),
    .X(_2594_));
 sky130_fd_sc_hd__inv_2 _5078_ (.A(_2594_),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _5079_ (.A(_2594_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _5080_ (.A(_2594_),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_2 _5081_ (.A(_2594_),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_2 _5082_ (.A(_2594_),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _5083_ (.A(_2594_),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_2 _5084_ (.A(_2594_),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_2 _5085_ (.A(_2594_),
    .Y(_0408_));
 sky130_fd_sc_hd__inv_2 _5086_ (.A(_2594_),
    .Y(_0409_));
 sky130_fd_sc_hd__inv_2 _5087_ (.A(_2594_),
    .Y(_0410_));
 sky130_fd_sc_hd__clkbuf_8 _5088_ (.A(_2591_),
    .X(_2595_));
 sky130_fd_sc_hd__inv_2 _5089_ (.A(_2595_),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_2 _5090_ (.A(_2595_),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_2 _5091_ (.A(_2595_),
    .Y(_0413_));
 sky130_fd_sc_hd__inv_2 _5092_ (.A(_2595_),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_2 _5093_ (.A(_2595_),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_2 _5094_ (.A(_2595_),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_2 _5095_ (.A(_2595_),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_2 _5096_ (.A(_2595_),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_2 _5097_ (.A(_2595_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _5098_ (.A(_2595_),
    .Y(_0420_));
 sky130_fd_sc_hd__buf_4 _5099_ (.A(_2591_),
    .X(_2596_));
 sky130_fd_sc_hd__inv_2 _5100_ (.A(_2596_),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _5101_ (.A(_2596_),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _5102_ (.A(_2596_),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _5103_ (.A(_2596_),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _5104_ (.A(_2596_),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _5105_ (.A(_2596_),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_2 _5106_ (.A(_2596_),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_2 _5107_ (.A(_2596_),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _5108_ (.A(_2596_),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _5109_ (.A(_2596_),
    .Y(_0430_));
 sky130_fd_sc_hd__clkbuf_8 _5110_ (.A(_2591_),
    .X(_2597_));
 sky130_fd_sc_hd__inv_2 _5111_ (.A(_2597_),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _5112_ (.A(_2597_),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _5113_ (.A(_2597_),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _5114_ (.A(_2597_),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _5115_ (.A(_2597_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _5116_ (.A(_2597_),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _5117_ (.A(_2597_),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _5118_ (.A(_2597_),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _5119_ (.A(_2597_),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _5120_ (.A(_2597_),
    .Y(_0440_));
 sky130_fd_sc_hd__clkbuf_8 _5121_ (.A(_2591_),
    .X(_2598_));
 sky130_fd_sc_hd__inv_2 _5122_ (.A(_2598_),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _5123_ (.A(_2598_),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_2 _5124_ (.A(_2598_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _5125_ (.A(_2598_),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _5126_ (.A(_2598_),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _5127_ (.A(_2598_),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_2 _5128_ (.A(_2598_),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_2 _5129_ (.A(_2598_),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_2 _5130_ (.A(_2598_),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_2 _5131_ (.A(_2598_),
    .Y(_0450_));
 sky130_fd_sc_hd__clkbuf_8 _5132_ (.A(_2591_),
    .X(_2599_));
 sky130_fd_sc_hd__inv_2 _5133_ (.A(_2599_),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _5134_ (.A(_2599_),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _5135_ (.A(_2599_),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _5136_ (.A(_2599_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _5137_ (.A(_2599_),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _5138_ (.A(_2599_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _5139_ (.A(_2599_),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _5140_ (.A(_2599_),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _5141_ (.A(_2599_),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _5142_ (.A(_2599_),
    .Y(_0460_));
 sky130_fd_sc_hd__clkbuf_8 _5143_ (.A(_2591_),
    .X(_2600_));
 sky130_fd_sc_hd__inv_2 _5144_ (.A(_2600_),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _5145_ (.A(_2600_),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _5146_ (.A(_2600_),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _5147_ (.A(_2600_),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _5148_ (.A(_2600_),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _5149_ (.A(_2600_),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _5150_ (.A(_2600_),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_2 _5151_ (.A(_2600_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _5152_ (.A(_2600_),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _5153_ (.A(_2600_),
    .Y(_0470_));
 sky130_fd_sc_hd__clkbuf_8 _5154_ (.A(_2591_),
    .X(_2601_));
 sky130_fd_sc_hd__inv_2 _5155_ (.A(_2601_),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _5156_ (.A(_2601_),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _5157_ (.A(_2601_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _5158_ (.A(_2601_),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_2 _5159_ (.A(_2601_),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _5160_ (.A(_2601_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _5161_ (.A(_2601_),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_2 _5162_ (.A(_2601_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _5163_ (.A(_2601_),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_2 _5164_ (.A(_2601_),
    .Y(_0480_));
 sky130_fd_sc_hd__clkbuf_8 _5165_ (.A(_2531_),
    .X(_2602_));
 sky130_fd_sc_hd__inv_2 _5166_ (.A(_2602_),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_2 _5167_ (.A(_2602_),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _5168_ (.A(_2602_),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _5169_ (.A(_2602_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _5170_ (.A(_2602_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _5171_ (.A(_2602_),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _5172_ (.A(_2602_),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_2 _5173_ (.A(_2602_),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _5174_ (.A(_2602_),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _5175_ (.A(_2602_),
    .Y(_0490_));
 sky130_fd_sc_hd__buf_4 _5176_ (.A(_2531_),
    .X(_2603_));
 sky130_fd_sc_hd__inv_2 _5177_ (.A(_2603_),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _5178_ (.A(_2603_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _5179_ (.A(_2603_),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _5180_ (.A(_2603_),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _5181_ (.A(_2603_),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _5182_ (.A(_2603_),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _5183_ (.A(_2603_),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _5184_ (.A(_2603_),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _5185_ (.A(_2603_),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _5186_ (.A(_2603_),
    .Y(_0500_));
 sky130_fd_sc_hd__clkbuf_8 _5187_ (.A(_2531_),
    .X(_2604_));
 sky130_fd_sc_hd__inv_2 _5188_ (.A(_2604_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _5189_ (.A(_2604_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _5190_ (.A(_2604_),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _5191_ (.A(_2604_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _5192_ (.A(_2604_),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _5193_ (.A(_2604_),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _5194_ (.A(_2604_),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _5195_ (.A(_2604_),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _5196_ (.A(_2604_),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _5197_ (.A(_2604_),
    .Y(_0510_));
 sky130_fd_sc_hd__buf_6 _5198_ (.A(_2531_),
    .X(_2605_));
 sky130_fd_sc_hd__inv_2 _5199_ (.A(_2605_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _5200_ (.A(_2605_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _5201_ (.A(_2605_),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _5202_ (.A(_2605_),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _5203_ (.A(_2605_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _5204_ (.A(_2605_),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _5205_ (.A(_2605_),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _5206_ (.A(_2605_),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _5207_ (.A(_2605_),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _5208_ (.A(_2605_),
    .Y(_0520_));
 sky130_fd_sc_hd__buf_6 _5209_ (.A(_2531_),
    .X(_2606_));
 sky130_fd_sc_hd__inv_2 _5210_ (.A(_2606_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _5211_ (.A(_2606_),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _5212_ (.A(_2606_),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _5213_ (.A(_2606_),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _5214_ (.A(_2606_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _5215_ (.A(_2606_),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _5216_ (.A(_2606_),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _5217_ (.A(_2606_),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _5218_ (.A(_2606_),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _5219_ (.A(_2606_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _5220_ (.A(_2549_),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _5221_ (.A(_2549_),
    .Y(_0532_));
 sky130_fd_sc_hd__dfxtp_2 _5222_ (.CLK(clknet_leaf_34_CLK),
    .D(_0533_),
    .Q(net19));
 sky130_fd_sc_hd__dfstp_1 _5223_ (.CLK(clknet_leaf_16_CLK),
    .D(_0534_),
    .SET_B(_0000_),
    .Q(\col_input[0] ));
 sky130_fd_sc_hd__dfrtp_2 _5224_ (.CLK(clknet_leaf_17_CLK),
    .D(_0535_),
    .RESET_B(_0001_),
    .Q(\col_input[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5225_ (.CLK(clknet_leaf_17_CLK),
    .D(_0536_),
    .RESET_B(_0002_),
    .Q(\col_input[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5226_ (.CLK(clknet_leaf_17_CLK),
    .D(_0537_),
    .RESET_B(_0003_),
    .Q(\col_input[3] ));
 sky130_fd_sc_hd__dfrtp_4 _5227_ (.CLK(clknet_leaf_17_CLK),
    .D(_0538_),
    .RESET_B(_0004_),
    .Q(\col_input[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5228_ (.CLK(clknet_leaf_21_CLK),
    .D(_0539_),
    .RESET_B(_0005_),
    .Q(\col_input[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5229_ (.CLK(clknet_leaf_18_CLK),
    .D(_0540_),
    .RESET_B(_0006_),
    .Q(\col_input[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5230_ (.CLK(clknet_leaf_18_CLK),
    .D(_0541_),
    .RESET_B(_0007_),
    .Q(\col_input[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5231_ (.CLK(clknet_leaf_20_CLK),
    .D(_0542_),
    .RESET_B(_0008_),
    .Q(\col_input[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5232_ (.CLK(clknet_leaf_21_CLK),
    .D(_0543_),
    .RESET_B(_0009_),
    .Q(\col_input[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5233_ (.CLK(clknet_leaf_20_CLK),
    .D(_0544_),
    .RESET_B(_0010_),
    .Q(\col_input[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5234_ (.CLK(clknet_leaf_20_CLK),
    .D(_0545_),
    .RESET_B(_0011_),
    .Q(\col_input[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5235_ (.CLK(clknet_leaf_21_CLK),
    .D(_0546_),
    .RESET_B(_0012_),
    .Q(\col_input[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5236_ (.CLK(clknet_leaf_21_CLK),
    .D(_0547_),
    .RESET_B(_0013_),
    .Q(\col_input[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5237_ (.CLK(clknet_leaf_21_CLK),
    .D(_0548_),
    .RESET_B(_0014_),
    .Q(\col_input[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5238_ (.CLK(clknet_leaf_21_CLK),
    .D(_0549_),
    .RESET_B(_0015_),
    .Q(\col_input[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5239_ (.CLK(clknet_leaf_21_CLK),
    .D(_0550_),
    .RESET_B(_0016_),
    .Q(\col_input[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5240_ (.CLK(clknet_leaf_21_CLK),
    .D(_0551_),
    .RESET_B(_0017_),
    .Q(\col_input[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5241_ (.CLK(clknet_leaf_21_CLK),
    .D(_0552_),
    .RESET_B(_0018_),
    .Q(\col_input[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5242_ (.CLK(clknet_leaf_21_CLK),
    .D(_0553_),
    .RESET_B(_0019_),
    .Q(\col_input[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5243_ (.CLK(clknet_leaf_22_CLK),
    .D(_0554_),
    .RESET_B(_0020_),
    .Q(\col_input[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5244_ (.CLK(clknet_leaf_22_CLK),
    .D(_0555_),
    .RESET_B(_0021_),
    .Q(\col_input[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5245_ (.CLK(clknet_leaf_22_CLK),
    .D(_0556_),
    .RESET_B(_0022_),
    .Q(\col_input[22] ));
 sky130_fd_sc_hd__dfrtp_1 _5246_ (.CLK(clknet_leaf_22_CLK),
    .D(_0557_),
    .RESET_B(_0023_),
    .Q(\col_input[23] ));
 sky130_fd_sc_hd__dfrtp_1 _5247_ (.CLK(clknet_leaf_22_CLK),
    .D(_0558_),
    .RESET_B(_0024_),
    .Q(\col_input[24] ));
 sky130_fd_sc_hd__dfrtp_1 _5248_ (.CLK(clknet_leaf_22_CLK),
    .D(_0559_),
    .RESET_B(_0025_),
    .Q(\col_input[25] ));
 sky130_fd_sc_hd__dfrtp_1 _5249_ (.CLK(clknet_leaf_22_CLK),
    .D(_0560_),
    .RESET_B(_0026_),
    .Q(\col_input[26] ));
 sky130_fd_sc_hd__dfrtp_1 _5250_ (.CLK(clknet_leaf_22_CLK),
    .D(_0561_),
    .RESET_B(_0027_),
    .Q(\col_input[27] ));
 sky130_fd_sc_hd__dfrtp_1 _5251_ (.CLK(clknet_leaf_22_CLK),
    .D(_0562_),
    .RESET_B(_0028_),
    .Q(\col_input[28] ));
 sky130_fd_sc_hd__dfrtp_1 _5252_ (.CLK(clknet_leaf_29_CLK),
    .D(_0563_),
    .RESET_B(_0029_),
    .Q(\col_input[29] ));
 sky130_fd_sc_hd__dfrtp_1 _5253_ (.CLK(clknet_leaf_29_CLK),
    .D(_0564_),
    .RESET_B(_0030_),
    .Q(\col_input[30] ));
 sky130_fd_sc_hd__dfrtp_1 _5254_ (.CLK(clknet_leaf_29_CLK),
    .D(_0565_),
    .RESET_B(_0031_),
    .Q(\col_input[31] ));
 sky130_fd_sc_hd__dfstp_1 _5255_ (.CLK(clknet_leaf_30_CLK),
    .D(_0566_),
    .SET_B(_0032_),
    .Q(\col_operation[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5256_ (.CLK(clknet_leaf_29_CLK),
    .D(_0567_),
    .RESET_B(_0033_),
    .Q(\col_operation[1] ));
 sky130_fd_sc_hd__dfrtp_2 _5257_ (.CLK(clknet_leaf_29_CLK),
    .D(_0568_),
    .RESET_B(_0034_),
    .Q(\col_operation[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5258_ (.CLK(clknet_leaf_29_CLK),
    .D(_0569_),
    .RESET_B(_0035_),
    .Q(\col_operation[3] ));
 sky130_fd_sc_hd__dfstp_4 _5259_ (.CLK(clknet_leaf_29_CLK),
    .D(_0570_),
    .SET_B(_0036_),
    .Q(\col_operation[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5260_ (.CLK(clknet_leaf_32_CLK),
    .D(_0571_),
    .RESET_B(_0037_),
    .Q(\valid_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5261_ (.CLK(clknet_leaf_32_CLK),
    .D(_0572_),
    .RESET_B(_0038_),
    .Q(\valid_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5262_ (.CLK(clknet_leaf_32_CLK),
    .D(_0573_),
    .RESET_B(_0039_),
    .Q(\valid_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5263_ (.CLK(clknet_leaf_32_CLK),
    .D(_0574_),
    .RESET_B(_0040_),
    .Q(\valid_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5264_ (.CLK(clknet_leaf_32_CLK),
    .D(_0575_),
    .RESET_B(_0041_),
    .Q(\valid_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5265_ (.CLK(clknet_leaf_32_CLK),
    .D(_0576_),
    .RESET_B(_0042_),
    .Q(\valid_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5266_ (.CLK(clknet_leaf_33_CLK),
    .D(_0577_),
    .RESET_B(_0043_),
    .Q(\valid_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5267_ (.CLK(clknet_leaf_32_CLK),
    .D(_0578_),
    .RESET_B(_0044_),
    .Q(\valid_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5268_ (.CLK(clknet_leaf_32_CLK),
    .D(_0579_),
    .RESET_B(_0045_),
    .Q(\valid_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5269_ (.CLK(clknet_leaf_33_CLK),
    .D(_0580_),
    .RESET_B(_0046_),
    .Q(\valid_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5270_ (.CLK(clknet_leaf_32_CLK),
    .D(_0581_),
    .RESET_B(_0047_),
    .Q(\valid_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5271_ (.CLK(clknet_leaf_32_CLK),
    .D(_0582_),
    .RESET_B(_0048_),
    .Q(\valid_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5272_ (.CLK(clknet_leaf_32_CLK),
    .D(_0583_),
    .RESET_B(_0049_),
    .Q(\valid_counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5273_ (.CLK(clknet_leaf_32_CLK),
    .D(_0584_),
    .RESET_B(_0050_),
    .Q(\valid_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5274_ (.CLK(clknet_leaf_33_CLK),
    .D(_0585_),
    .RESET_B(_0051_),
    .Q(\valid_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5275_ (.CLK(clknet_leaf_33_CLK),
    .D(_0586_),
    .RESET_B(_0052_),
    .Q(\valid_counter[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5276_ (.CLK(clknet_leaf_33_CLK),
    .D(_0587_),
    .RESET_B(_0053_),
    .Q(\valid_counter[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5277_ (.CLK(clknet_leaf_33_CLK),
    .D(_0588_),
    .RESET_B(_0054_),
    .Q(\valid_counter[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5278_ (.CLK(clknet_leaf_33_CLK),
    .D(_0589_),
    .RESET_B(_0055_),
    .Q(\valid_counter[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5279_ (.CLK(clknet_leaf_33_CLK),
    .D(_0590_),
    .RESET_B(_0056_),
    .Q(\valid_counter[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5280_ (.CLK(clknet_leaf_33_CLK),
    .D(_0591_),
    .RESET_B(_0057_),
    .Q(\valid_counter[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5281_ (.CLK(clknet_leaf_33_CLK),
    .D(_0592_),
    .RESET_B(_0058_),
    .Q(\valid_counter[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5282_ (.CLK(clknet_leaf_33_CLK),
    .D(_0593_),
    .RESET_B(_0059_),
    .Q(\valid_counter[22] ));
 sky130_fd_sc_hd__dfrtp_1 _5283_ (.CLK(clknet_leaf_33_CLK),
    .D(_0594_),
    .RESET_B(_0060_),
    .Q(\valid_counter[23] ));
 sky130_fd_sc_hd__dfrtp_1 _5284_ (.CLK(clknet_leaf_34_CLK),
    .D(_0595_),
    .RESET_B(_0061_),
    .Q(\valid_counter[24] ));
 sky130_fd_sc_hd__dfrtp_1 _5285_ (.CLK(clknet_leaf_33_CLK),
    .D(_0596_),
    .RESET_B(_0062_),
    .Q(\valid_counter[25] ));
 sky130_fd_sc_hd__dfrtp_1 _5286_ (.CLK(clknet_leaf_33_CLK),
    .D(_0597_),
    .RESET_B(_0063_),
    .Q(\valid_counter[26] ));
 sky130_fd_sc_hd__dfrtp_1 _5287_ (.CLK(clknet_leaf_34_CLK),
    .D(_0598_),
    .RESET_B(_0064_),
    .Q(\valid_counter[27] ));
 sky130_fd_sc_hd__dfrtp_1 _5288_ (.CLK(clknet_leaf_34_CLK),
    .D(_0599_),
    .RESET_B(_0065_),
    .Q(\valid_counter[28] ));
 sky130_fd_sc_hd__dfrtp_1 _5289_ (.CLK(clknet_leaf_34_CLK),
    .D(_0600_),
    .RESET_B(_0066_),
    .Q(\valid_counter[29] ));
 sky130_fd_sc_hd__dfrtp_1 _5290_ (.CLK(clknet_leaf_34_CLK),
    .D(_0601_),
    .RESET_B(_0067_),
    .Q(\valid_counter[30] ));
 sky130_fd_sc_hd__dfrtp_1 _5291_ (.CLK(clknet_leaf_34_CLK),
    .D(_0602_),
    .RESET_B(_0068_),
    .Q(\valid_counter[31] ));
 sky130_fd_sc_hd__dfrtp_1 _5292_ (.CLK(clknet_leaf_34_CLK),
    .D(_0603_),
    .RESET_B(_0069_),
    .Q(\k[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5293_ (.CLK(clknet_leaf_34_CLK),
    .D(_0604_),
    .RESET_B(_0070_),
    .Q(\k[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5294_ (.CLK(clknet_leaf_34_CLK),
    .D(_0605_),
    .RESET_B(_0071_),
    .Q(\k[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5295_ (.CLK(clknet_leaf_34_CLK),
    .D(_0606_),
    .RESET_B(_0072_),
    .Q(\k[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5296_ (.CLK(clknet_leaf_34_CLK),
    .D(_0607_),
    .RESET_B(_0073_),
    .Q(\k[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5297_ (.CLK(clknet_leaf_36_CLK),
    .D(_0608_),
    .RESET_B(_0074_),
    .Q(\k[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5298_ (.CLK(clknet_leaf_36_CLK),
    .D(_0609_),
    .RESET_B(_0075_),
    .Q(\k[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5299_ (.CLK(clknet_leaf_36_CLK),
    .D(_0610_),
    .RESET_B(_0076_),
    .Q(\k[7] ));
 sky130_fd_sc_hd__dfrtp_1 _5300_ (.CLK(clknet_leaf_38_CLK),
    .D(_0611_),
    .RESET_B(_0077_),
    .Q(\k[8] ));
 sky130_fd_sc_hd__dfrtp_1 _5301_ (.CLK(clknet_leaf_38_CLK),
    .D(_0612_),
    .RESET_B(_0078_),
    .Q(\k[9] ));
 sky130_fd_sc_hd__dfrtp_1 _5302_ (.CLK(clknet_leaf_38_CLK),
    .D(_0613_),
    .RESET_B(_0079_),
    .Q(\k[10] ));
 sky130_fd_sc_hd__dfrtp_1 _5303_ (.CLK(clknet_leaf_38_CLK),
    .D(_0614_),
    .RESET_B(_0080_),
    .Q(\k[11] ));
 sky130_fd_sc_hd__dfrtp_1 _5304_ (.CLK(clknet_leaf_38_CLK),
    .D(_0615_),
    .RESET_B(_0081_),
    .Q(\k[12] ));
 sky130_fd_sc_hd__dfrtp_1 _5305_ (.CLK(clknet_leaf_38_CLK),
    .D(_0616_),
    .RESET_B(_0082_),
    .Q(\k[13] ));
 sky130_fd_sc_hd__dfrtp_1 _5306_ (.CLK(clknet_leaf_38_CLK),
    .D(_0617_),
    .RESET_B(_0083_),
    .Q(\k[14] ));
 sky130_fd_sc_hd__dfrtp_1 _5307_ (.CLK(clknet_leaf_38_CLK),
    .D(_0618_),
    .RESET_B(_0084_),
    .Q(\k[15] ));
 sky130_fd_sc_hd__dfrtp_1 _5308_ (.CLK(clknet_leaf_38_CLK),
    .D(_0619_),
    .RESET_B(_0085_),
    .Q(\k[16] ));
 sky130_fd_sc_hd__dfrtp_1 _5309_ (.CLK(clknet_leaf_38_CLK),
    .D(_0620_),
    .RESET_B(_0086_),
    .Q(\k[17] ));
 sky130_fd_sc_hd__dfrtp_1 _5310_ (.CLK(clknet_leaf_38_CLK),
    .D(_0621_),
    .RESET_B(_0087_),
    .Q(\k[18] ));
 sky130_fd_sc_hd__dfrtp_1 _5311_ (.CLK(clknet_leaf_38_CLK),
    .D(_0622_),
    .RESET_B(_0088_),
    .Q(\k[19] ));
 sky130_fd_sc_hd__dfrtp_1 _5312_ (.CLK(clknet_leaf_38_CLK),
    .D(_0623_),
    .RESET_B(_0089_),
    .Q(\k[20] ));
 sky130_fd_sc_hd__dfrtp_1 _5313_ (.CLK(clknet_leaf_38_CLK),
    .D(_0624_),
    .RESET_B(_0090_),
    .Q(\k[21] ));
 sky130_fd_sc_hd__dfrtp_1 _5314_ (.CLK(clknet_leaf_38_CLK),
    .D(_0625_),
    .RESET_B(_0091_),
    .Q(\k[22] ));
 sky130_fd_sc_hd__dfrtp_1 _5315_ (.CLK(clknet_leaf_37_CLK),
    .D(_0626_),
    .RESET_B(_0092_),
    .Q(\k[23] ));
 sky130_fd_sc_hd__dfrtp_1 _5316_ (.CLK(clknet_leaf_37_CLK),
    .D(_0627_),
    .RESET_B(_0093_),
    .Q(\k[24] ));
 sky130_fd_sc_hd__dfrtp_1 _5317_ (.CLK(clknet_leaf_37_CLK),
    .D(_0628_),
    .RESET_B(_0094_),
    .Q(\k[25] ));
 sky130_fd_sc_hd__dfrtp_1 _5318_ (.CLK(clknet_leaf_37_CLK),
    .D(_0629_),
    .RESET_B(_0095_),
    .Q(\k[26] ));
 sky130_fd_sc_hd__dfrtp_1 _5319_ (.CLK(clknet_leaf_37_CLK),
    .D(_0630_),
    .RESET_B(_0096_),
    .Q(\k[27] ));
 sky130_fd_sc_hd__dfrtp_1 _5320_ (.CLK(clknet_leaf_36_CLK),
    .D(_0631_),
    .RESET_B(_0097_),
    .Q(\k[28] ));
 sky130_fd_sc_hd__dfrtp_1 _5321_ (.CLK(clknet_leaf_37_CLK),
    .D(_0632_),
    .RESET_B(_0098_),
    .Q(\k[29] ));
 sky130_fd_sc_hd__dfrtp_1 _5322_ (.CLK(clknet_leaf_37_CLK),
    .D(_0633_),
    .RESET_B(_0099_),
    .Q(\k[30] ));
 sky130_fd_sc_hd__dfrtp_1 _5323_ (.CLK(clknet_leaf_37_CLK),
    .D(_0634_),
    .RESET_B(_0100_),
    .Q(\k[31] ));
 sky130_fd_sc_hd__dfrtp_1 _5324_ (.CLK(clknet_leaf_20_CLK),
    .D(_0635_),
    .RESET_B(_0101_),
    .Q(\first_row[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5325_ (.CLK(clknet_leaf_20_CLK),
    .D(_0636_),
    .RESET_B(_0102_),
    .Q(\first_row[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5326_ (.CLK(clknet_leaf_24_CLK),
    .D(_0637_),
    .RESET_B(_0103_),
    .Q(\first_row[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5327_ (.CLK(clknet_leaf_7_CLK),
    .D(_0638_),
    .RESET_B(_0104_),
    .Q(\first_row[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5328_ (.CLK(clknet_leaf_3_CLK),
    .D(_0639_),
    .RESET_B(_0105_),
    .Q(\first_row[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5329_ (.CLK(clknet_leaf_8_CLK),
    .D(_0640_),
    .RESET_B(_0106_),
    .Q(\first_row[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5330_ (.CLK(clknet_leaf_3_CLK),
    .D(_0641_),
    .RESET_B(_0107_),
    .Q(\first_row[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5331_ (.CLK(clknet_leaf_6_CLK),
    .D(_0642_),
    .RESET_B(_0108_),
    .Q(\first_row[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5332_ (.CLK(clknet_leaf_20_CLK),
    .D(_0643_),
    .RESET_B(_0109_),
    .Q(\first_row[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5333_ (.CLK(clknet_leaf_20_CLK),
    .D(_0644_),
    .RESET_B(_0110_),
    .Q(\first_row[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5334_ (.CLK(clknet_leaf_24_CLK),
    .D(_0645_),
    .RESET_B(_0111_),
    .Q(\first_row[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5335_ (.CLK(clknet_leaf_7_CLK),
    .D(_0646_),
    .RESET_B(_0112_),
    .Q(\first_row[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5336_ (.CLK(clknet_leaf_7_CLK),
    .D(_0647_),
    .RESET_B(_0113_),
    .Q(\first_row[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5337_ (.CLK(clknet_leaf_10_CLK),
    .D(_0648_),
    .RESET_B(_0114_),
    .Q(\first_row[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5338_ (.CLK(clknet_leaf_6_CLK),
    .D(_0649_),
    .RESET_B(_0115_),
    .Q(\first_row[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5339_ (.CLK(clknet_leaf_7_CLK),
    .D(_0650_),
    .RESET_B(_0116_),
    .Q(\first_row[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5340_ (.CLK(clknet_leaf_22_CLK),
    .D(_0651_),
    .RESET_B(_0117_),
    .Q(\first_row[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5341_ (.CLK(clknet_leaf_22_CLK),
    .D(_0652_),
    .RESET_B(_0118_),
    .Q(\first_row[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5342_ (.CLK(clknet_leaf_25_CLK),
    .D(_0653_),
    .RESET_B(_0119_),
    .Q(\first_row[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5343_ (.CLK(clknet_leaf_7_CLK),
    .D(_0654_),
    .RESET_B(_0120_),
    .Q(\first_row[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5344_ (.CLK(clknet_leaf_5_CLK),
    .D(_0655_),
    .RESET_B(_0121_),
    .Q(\first_row[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5345_ (.CLK(clknet_leaf_6_CLK),
    .D(_0656_),
    .RESET_B(_0122_),
    .Q(\first_row[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5346_ (.CLK(clknet_leaf_5_CLK),
    .D(_0657_),
    .RESET_B(_0123_),
    .Q(\first_row[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5347_ (.CLK(clknet_leaf_6_CLK),
    .D(_0658_),
    .RESET_B(_0124_),
    .Q(\first_row[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5348_ (.CLK(clknet_leaf_28_CLK),
    .D(_0659_),
    .RESET_B(_0125_),
    .Q(\first_row[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5349_ (.CLK(clknet_leaf_31_CLK),
    .D(_0660_),
    .RESET_B(_0126_),
    .Q(\first_row[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5350_ (.CLK(clknet_leaf_23_CLK),
    .D(_0661_),
    .RESET_B(_0127_),
    .Q(\first_row[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5351_ (.CLK(clknet_leaf_7_CLK),
    .D(_0662_),
    .RESET_B(_0128_),
    .Q(\first_row[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5352_ (.CLK(clknet_leaf_43_CLK),
    .D(_0663_),
    .RESET_B(_0129_),
    .Q(\first_row[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5353_ (.CLK(clknet_leaf_44_CLK),
    .D(_0664_),
    .RESET_B(_0130_),
    .Q(\first_row[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5354_ (.CLK(clknet_leaf_47_CLK),
    .D(_0665_),
    .RESET_B(_0131_),
    .Q(\first_row[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5355_ (.CLK(clknet_leaf_47_CLK),
    .D(_0666_),
    .RESET_B(_0132_),
    .Q(\first_row[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5356_ (.CLK(clknet_leaf_31_CLK),
    .D(_0667_),
    .RESET_B(_0133_),
    .Q(\first_row[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5357_ (.CLK(clknet_leaf_35_CLK),
    .D(_0668_),
    .RESET_B(_0134_),
    .Q(\first_row[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5358_ (.CLK(clknet_leaf_35_CLK),
    .D(_0669_),
    .RESET_B(_0135_),
    .Q(\first_row[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5359_ (.CLK(clknet_leaf_39_CLK),
    .D(_0670_),
    .RESET_B(_0136_),
    .Q(\first_row[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5360_ (.CLK(clknet_leaf_44_CLK),
    .D(_0671_),
    .RESET_B(_0137_),
    .Q(\first_row[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5361_ (.CLK(clknet_leaf_47_CLK),
    .D(_0672_),
    .RESET_B(_0138_),
    .Q(\first_row[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5362_ (.CLK(clknet_leaf_47_CLK),
    .D(_0673_),
    .RESET_B(_0139_),
    .Q(\first_row[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5363_ (.CLK(clknet_leaf_47_CLK),
    .D(_0674_),
    .RESET_B(_0140_),
    .Q(\first_row[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5364_ (.CLK(clknet_leaf_31_CLK),
    .D(_0675_),
    .RESET_B(_0141_),
    .Q(\first_row[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5365_ (.CLK(clknet_leaf_31_CLK),
    .D(_0676_),
    .RESET_B(_0142_),
    .Q(\first_row[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5366_ (.CLK(clknet_leaf_35_CLK),
    .D(_0677_),
    .RESET_B(_0143_),
    .Q(\first_row[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5367_ (.CLK(clknet_leaf_40_CLK),
    .D(_0678_),
    .RESET_B(_0144_),
    .Q(\first_row[6][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5368_ (.CLK(clknet_leaf_44_CLK),
    .D(_0679_),
    .RESET_B(_0145_),
    .Q(\first_row[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5369_ (.CLK(clknet_leaf_47_CLK),
    .D(_0680_),
    .RESET_B(_0146_),
    .Q(\first_row[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5370_ (.CLK(clknet_leaf_47_CLK),
    .D(_0681_),
    .RESET_B(_0147_),
    .Q(\first_row[6][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5371_ (.CLK(clknet_leaf_44_CLK),
    .D(_0682_),
    .RESET_B(_0148_),
    .Q(\first_row[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5372_ (.CLK(clknet_leaf_30_CLK),
    .D(_0683_),
    .RESET_B(_0149_),
    .Q(\first_row[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5373_ (.CLK(clknet_leaf_29_CLK),
    .D(_0684_),
    .RESET_B(_0150_),
    .Q(\first_row[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5374_ (.CLK(clknet_leaf_8_CLK),
    .D(_0685_),
    .RESET_B(_0151_),
    .Q(\first_row[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5375_ (.CLK(clknet_leaf_20_CLK),
    .D(_0686_),
    .RESET_B(_0152_),
    .Q(\first_row[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5376_ (.CLK(clknet_leaf_20_CLK),
    .D(_0687_),
    .RESET_B(_0153_),
    .Q(\first_row[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5377_ (.CLK(clknet_leaf_8_CLK),
    .D(_0688_),
    .RESET_B(_0154_),
    .Q(\first_row[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5378_ (.CLK(clknet_leaf_8_CLK),
    .D(_0689_),
    .RESET_B(_0155_),
    .Q(\first_row[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5379_ (.CLK(clknet_leaf_8_CLK),
    .D(_0690_),
    .RESET_B(_0156_),
    .Q(\first_row[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5380_ (.CLK(clknet_leaf_18_CLK),
    .D(_0691_),
    .RESET_B(_0157_),
    .Q(\first_row[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5381_ (.CLK(clknet_leaf_18_CLK),
    .D(_0692_),
    .RESET_B(_0158_),
    .Q(\first_row[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5382_ (.CLK(clknet_leaf_8_CLK),
    .D(_0693_),
    .RESET_B(_0159_),
    .Q(\first_row[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5383_ (.CLK(clknet_leaf_8_CLK),
    .D(_0694_),
    .RESET_B(_0160_),
    .Q(\first_row[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5384_ (.CLK(clknet_leaf_1_CLK),
    .D(_0695_),
    .RESET_B(_0161_),
    .Q(\first_row[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5385_ (.CLK(clknet_leaf_62_CLK),
    .D(_0696_),
    .RESET_B(_0162_),
    .Q(\first_row[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5386_ (.CLK(clknet_leaf_63_CLK),
    .D(_0697_),
    .RESET_B(_0163_),
    .Q(\first_row[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5387_ (.CLK(clknet_leaf_63_CLK),
    .D(_0698_),
    .RESET_B(_0164_),
    .Q(\first_row[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5388_ (.CLK(clknet_leaf_19_CLK),
    .D(_0699_),
    .RESET_B(_0165_),
    .Q(\first_row[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5389_ (.CLK(clknet_leaf_13_CLK),
    .D(_0700_),
    .RESET_B(_0166_),
    .Q(\first_row[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5390_ (.CLK(clknet_leaf_13_CLK),
    .D(_0701_),
    .RESET_B(_0167_),
    .Q(\first_row[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5391_ (.CLK(clknet_leaf_9_CLK),
    .D(_0702_),
    .RESET_B(_0168_),
    .Q(\first_row[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5392_ (.CLK(clknet_leaf_1_CLK),
    .D(_0703_),
    .RESET_B(_0169_),
    .Q(\first_row[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5393_ (.CLK(clknet_leaf_63_CLK),
    .D(_0704_),
    .RESET_B(_0170_),
    .Q(\first_row[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5394_ (.CLK(clknet_leaf_62_CLK),
    .D(_0705_),
    .RESET_B(_0171_),
    .Q(\first_row[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5395_ (.CLK(clknet_leaf_62_CLK),
    .D(_0706_),
    .RESET_B(_0172_),
    .Q(\first_row[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5396_ (.CLK(clknet_leaf_13_CLK),
    .D(_0707_),
    .RESET_B(_0173_),
    .Q(\first_row[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5397_ (.CLK(clknet_leaf_20_CLK),
    .D(_0708_),
    .RESET_B(_0174_),
    .Q(\first_row[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5398_ (.CLK(clknet_leaf_13_CLK),
    .D(_0709_),
    .RESET_B(_0175_),
    .Q(\first_row[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5399_ (.CLK(clknet_leaf_10_CLK),
    .D(_0710_),
    .RESET_B(_0176_),
    .Q(\first_row[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5400_ (.CLK(clknet_leaf_1_CLK),
    .D(_0711_),
    .RESET_B(_0177_),
    .Q(\first_row[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5401_ (.CLK(clknet_leaf_62_CLK),
    .D(_0712_),
    .RESET_B(_0178_),
    .Q(\first_row[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5402_ (.CLK(clknet_leaf_62_CLK),
    .D(_0713_),
    .RESET_B(_0179_),
    .Q(\first_row[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5403_ (.CLK(clknet_leaf_62_CLK),
    .D(_0714_),
    .RESET_B(_0180_),
    .Q(\first_row[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5404_ (.CLK(clknet_leaf_16_CLK),
    .D(_0715_),
    .RESET_B(_0181_),
    .Q(\first_row[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5405_ (.CLK(clknet_leaf_16_CLK),
    .D(_0716_),
    .RESET_B(_0182_),
    .Q(\first_row[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5406_ (.CLK(clknet_leaf_14_CLK),
    .D(_0717_),
    .RESET_B(_0183_),
    .Q(\first_row[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5407_ (.CLK(clknet_leaf_11_CLK),
    .D(_0718_),
    .RESET_B(_0184_),
    .Q(\first_row[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5408_ (.CLK(clknet_leaf_2_CLK),
    .D(_0719_),
    .RESET_B(_0185_),
    .Q(\first_row[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5409_ (.CLK(clknet_leaf_11_CLK),
    .D(_0720_),
    .RESET_B(_0186_),
    .Q(\first_row[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5410_ (.CLK(clknet_leaf_3_CLK),
    .D(_0721_),
    .RESET_B(_0187_),
    .Q(\first_row[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5411_ (.CLK(clknet_leaf_2_CLK),
    .D(_0722_),
    .RESET_B(_0188_),
    .Q(\first_row[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5412_ (.CLK(clknet_leaf_16_CLK),
    .D(_0723_),
    .RESET_B(_0189_),
    .Q(\first_row[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5413_ (.CLK(clknet_leaf_16_CLK),
    .D(_0724_),
    .RESET_B(_0190_),
    .Q(\first_row[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5414_ (.CLK(clknet_leaf_14_CLK),
    .D(_0725_),
    .RESET_B(_0191_),
    .Q(\first_row[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5415_ (.CLK(clknet_leaf_11_CLK),
    .D(_0726_),
    .RESET_B(_0192_),
    .Q(\first_row[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5416_ (.CLK(clknet_leaf_1_CLK),
    .D(_0727_),
    .RESET_B(_0193_),
    .Q(\first_row[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5417_ (.CLK(clknet_leaf_63_CLK),
    .D(_0728_),
    .RESET_B(_0194_),
    .Q(\first_row[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5418_ (.CLK(clknet_leaf_63_CLK),
    .D(_0729_),
    .RESET_B(_0195_),
    .Q(\first_row[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5419_ (.CLK(clknet_leaf_63_CLK),
    .D(_0730_),
    .RESET_B(_0196_),
    .Q(\first_row[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5420_ (.CLK(clknet_leaf_13_CLK),
    .D(_0731_),
    .RESET_B(_0197_),
    .Q(\first_row[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5421_ (.CLK(clknet_leaf_19_CLK),
    .D(_0732_),
    .RESET_B(_0198_),
    .Q(\first_row[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5422_ (.CLK(clknet_leaf_13_CLK),
    .D(_0733_),
    .RESET_B(_0199_),
    .Q(\first_row[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5423_ (.CLK(clknet_leaf_10_CLK),
    .D(_0734_),
    .RESET_B(_0200_),
    .Q(\first_row[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5424_ (.CLK(clknet_leaf_1_CLK),
    .D(_0735_),
    .RESET_B(_0201_),
    .Q(\first_row[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5425_ (.CLK(clknet_leaf_62_CLK),
    .D(_0736_),
    .RESET_B(_0202_),
    .Q(\first_row[13][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5426_ (.CLK(clknet_leaf_0_CLK),
    .D(_0737_),
    .RESET_B(_0203_),
    .Q(\first_row[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5427_ (.CLK(clknet_leaf_62_CLK),
    .D(_0738_),
    .RESET_B(_0204_),
    .Q(\first_row[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5428_ (.CLK(clknet_leaf_19_CLK),
    .D(_0739_),
    .RESET_B(_0205_),
    .Q(\first_row[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5429_ (.CLK(clknet_leaf_19_CLK),
    .D(_0740_),
    .RESET_B(_0206_),
    .Q(\first_row[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5430_ (.CLK(clknet_leaf_13_CLK),
    .D(_0741_),
    .RESET_B(_0207_),
    .Q(\first_row[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5431_ (.CLK(clknet_leaf_8_CLK),
    .D(_0742_),
    .RESET_B(_0208_),
    .Q(\first_row[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5432_ (.CLK(clknet_leaf_1_CLK),
    .D(_0743_),
    .RESET_B(_0209_),
    .Q(\first_row[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5433_ (.CLK(clknet_leaf_1_CLK),
    .D(_0744_),
    .RESET_B(_0210_),
    .Q(\first_row[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5434_ (.CLK(clknet_leaf_0_CLK),
    .D(_0745_),
    .RESET_B(_0211_),
    .Q(\first_row[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5435_ (.CLK(clknet_leaf_0_CLK),
    .D(_0746_),
    .RESET_B(_0212_),
    .Q(\first_row[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5436_ (.CLK(clknet_leaf_19_CLK),
    .D(_0747_),
    .RESET_B(_0213_),
    .Q(\first_row[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5437_ (.CLK(clknet_leaf_19_CLK),
    .D(_0748_),
    .RESET_B(_0214_),
    .Q(\first_row[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5438_ (.CLK(clknet_leaf_13_CLK),
    .D(_0749_),
    .RESET_B(_0215_),
    .Q(\first_row[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5439_ (.CLK(clknet_leaf_9_CLK),
    .D(_0750_),
    .RESET_B(_0216_),
    .Q(\first_row[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5440_ (.CLK(clknet_leaf_3_CLK),
    .D(_0751_),
    .RESET_B(_0217_),
    .Q(\first_row[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5441_ (.CLK(clknet_leaf_9_CLK),
    .D(_0752_),
    .RESET_B(_0218_),
    .Q(\first_row[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5442_ (.CLK(clknet_leaf_3_CLK),
    .D(_0753_),
    .RESET_B(_0219_),
    .Q(\first_row[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5443_ (.CLK(clknet_leaf_3_CLK),
    .D(_0754_),
    .RESET_B(_0220_),
    .Q(\first_row[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5444_ (.CLK(clknet_leaf_16_CLK),
    .D(_0755_),
    .RESET_B(_0221_),
    .Q(\first_row[16][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5445_ (.CLK(clknet_leaf_16_CLK),
    .D(_0756_),
    .RESET_B(_0222_),
    .Q(\first_row[16][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5446_ (.CLK(clknet_leaf_17_CLK),
    .D(_0757_),
    .RESET_B(_0223_),
    .Q(\first_row[16][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5447_ (.CLK(clknet_leaf_16_CLK),
    .D(_0758_),
    .RESET_B(_0224_),
    .Q(\first_row[16][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5448_ (.CLK(clknet_leaf_16_CLK),
    .D(_0759_),
    .RESET_B(_0225_),
    .Q(\first_row[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5449_ (.CLK(clknet_leaf_17_CLK),
    .D(_0760_),
    .RESET_B(_0226_),
    .Q(\first_row[16][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5450_ (.CLK(clknet_leaf_17_CLK),
    .D(_0761_),
    .RESET_B(_0227_),
    .Q(\first_row[16][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5451_ (.CLK(clknet_leaf_17_CLK),
    .D(_0762_),
    .RESET_B(_0228_),
    .Q(\first_row[16][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5452_ (.CLK(clknet_leaf_13_CLK),
    .D(_0763_),
    .RESET_B(_0229_),
    .Q(\first_row[17][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5453_ (.CLK(clknet_leaf_17_CLK),
    .D(_0764_),
    .RESET_B(_0230_),
    .Q(\first_row[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5454_ (.CLK(clknet_leaf_12_CLK),
    .D(_0765_),
    .RESET_B(_0231_),
    .Q(\first_row[17][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5455_ (.CLK(clknet_leaf_10_CLK),
    .D(_0766_),
    .RESET_B(_0232_),
    .Q(\first_row[17][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5456_ (.CLK(clknet_leaf_1_CLK),
    .D(_0767_),
    .RESET_B(_0233_),
    .Q(\first_row[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5457_ (.CLK(clknet_leaf_4_CLK),
    .D(_0768_),
    .RESET_B(_0234_),
    .Q(\first_row[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5458_ (.CLK(clknet_leaf_1_CLK),
    .D(_0769_),
    .RESET_B(_0235_),
    .Q(\first_row[17][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5459_ (.CLK(clknet_leaf_4_CLK),
    .D(_0770_),
    .RESET_B(_0236_),
    .Q(\first_row[17][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5460_ (.CLK(clknet_leaf_15_CLK),
    .D(_0771_),
    .RESET_B(_0237_),
    .Q(\second_row[0][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5461_ (.CLK(clknet_leaf_15_CLK),
    .D(_0772_),
    .RESET_B(_0238_),
    .Q(\second_row[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5462_ (.CLK(clknet_leaf_12_CLK),
    .D(_0773_),
    .RESET_B(_0239_),
    .Q(\second_row[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5463_ (.CLK(clknet_leaf_11_CLK),
    .D(_0774_),
    .RESET_B(_0240_),
    .Q(\second_row[0][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5464_ (.CLK(clknet_leaf_2_CLK),
    .D(_0775_),
    .RESET_B(_0241_),
    .Q(\second_row[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5465_ (.CLK(clknet_leaf_64_CLK),
    .D(_0776_),
    .RESET_B(_0242_),
    .Q(\second_row[0][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5466_ (.CLK(clknet_leaf_0_CLK),
    .D(_0777_),
    .RESET_B(_0243_),
    .Q(\second_row[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5467_ (.CLK(clknet_leaf_64_CLK),
    .D(_0778_),
    .RESET_B(_0244_),
    .Q(\second_row[0][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5468_ (.CLK(clknet_leaf_23_CLK),
    .D(_0779_),
    .RESET_B(_0245_),
    .Q(\second_row[1][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5469_ (.CLK(clknet_leaf_23_CLK),
    .D(_0780_),
    .RESET_B(_0246_),
    .Q(\second_row[1][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5470_ (.CLK(clknet_leaf_24_CLK),
    .D(_0781_),
    .RESET_B(_0247_),
    .Q(\second_row[1][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5471_ (.CLK(clknet_leaf_7_CLK),
    .D(_0782_),
    .RESET_B(_0248_),
    .Q(\second_row[1][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5472_ (.CLK(clknet_leaf_3_CLK),
    .D(_0783_),
    .RESET_B(_0249_),
    .Q(\second_row[1][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5473_ (.CLK(clknet_leaf_9_CLK),
    .D(_0784_),
    .RESET_B(_0250_),
    .Q(\second_row[1][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5474_ (.CLK(clknet_leaf_3_CLK),
    .D(_0785_),
    .RESET_B(_0251_),
    .Q(\second_row[1][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5475_ (.CLK(clknet_leaf_5_CLK),
    .D(_0786_),
    .RESET_B(_0252_),
    .Q(\second_row[1][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5476_ (.CLK(clknet_leaf_23_CLK),
    .D(_0787_),
    .RESET_B(_0253_),
    .Q(\second_row[2][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5477_ (.CLK(clknet_leaf_23_CLK),
    .D(_0788_),
    .RESET_B(_0254_),
    .Q(\second_row[2][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5478_ (.CLK(clknet_leaf_24_CLK),
    .D(_0789_),
    .RESET_B(_0255_),
    .Q(\second_row[2][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5479_ (.CLK(clknet_leaf_7_CLK),
    .D(_0790_),
    .RESET_B(_0256_),
    .Q(\second_row[2][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5480_ (.CLK(clknet_leaf_24_CLK),
    .D(_0791_),
    .RESET_B(_0257_),
    .Q(\second_row[2][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5481_ (.CLK(clknet_leaf_6_CLK),
    .D(_0792_),
    .RESET_B(_0258_),
    .Q(\second_row[2][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5482_ (.CLK(clknet_leaf_6_CLK),
    .D(_0793_),
    .RESET_B(_0259_),
    .Q(\second_row[2][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5483_ (.CLK(clknet_leaf_6_CLK),
    .D(_0794_),
    .RESET_B(_0260_),
    .Q(\second_row[2][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5484_ (.CLK(clknet_leaf_28_CLK),
    .D(_0795_),
    .RESET_B(_0261_),
    .Q(\second_row[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5485_ (.CLK(clknet_leaf_22_CLK),
    .D(_0796_),
    .RESET_B(_0262_),
    .Q(\second_row[3][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5486_ (.CLK(clknet_leaf_25_CLK),
    .D(_0797_),
    .RESET_B(_0263_),
    .Q(\second_row[3][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5487_ (.CLK(clknet_leaf_7_CLK),
    .D(_0798_),
    .RESET_B(_0264_),
    .Q(\second_row[3][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5488_ (.CLK(clknet_leaf_6_CLK),
    .D(_0799_),
    .RESET_B(_0265_),
    .Q(\second_row[3][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5489_ (.CLK(clknet_leaf_57_CLK),
    .D(_0800_),
    .RESET_B(_0266_),
    .Q(\second_row[3][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5490_ (.CLK(clknet_leaf_6_CLK),
    .D(_0801_),
    .RESET_B(_0267_),
    .Q(\second_row[3][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5491_ (.CLK(clknet_leaf_57_CLK),
    .D(_0802_),
    .RESET_B(_0268_),
    .Q(\second_row[3][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5492_ (.CLK(clknet_leaf_28_CLK),
    .D(_0803_),
    .RESET_B(_0269_),
    .Q(\second_row[4][0] ));
 sky130_fd_sc_hd__dfrtp_2 _5493_ (.CLK(clknet_leaf_31_CLK),
    .D(_0804_),
    .RESET_B(_0270_),
    .Q(\second_row[4][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5494_ (.CLK(clknet_leaf_25_CLK),
    .D(_0805_),
    .RESET_B(_0271_),
    .Q(\second_row[4][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5495_ (.CLK(clknet_leaf_7_CLK),
    .D(_0806_),
    .RESET_B(_0272_),
    .Q(\second_row[4][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5496_ (.CLK(clknet_leaf_44_CLK),
    .D(_0807_),
    .RESET_B(_0273_),
    .Q(\second_row[4][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5497_ (.CLK(clknet_leaf_44_CLK),
    .D(_0808_),
    .RESET_B(_0274_),
    .Q(\second_row[4][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5498_ (.CLK(clknet_leaf_47_CLK),
    .D(_0809_),
    .RESET_B(_0275_),
    .Q(\second_row[4][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5499_ (.CLK(clknet_leaf_49_CLK),
    .D(_0810_),
    .RESET_B(_0276_),
    .Q(\second_row[4][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5500_ (.CLK(clknet_leaf_35_CLK),
    .D(_0811_),
    .RESET_B(_0277_),
    .Q(\second_row[5][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5501_ (.CLK(clknet_leaf_35_CLK),
    .D(_0812_),
    .RESET_B(_0278_),
    .Q(\second_row[5][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5502_ (.CLK(clknet_leaf_35_CLK),
    .D(_0813_),
    .RESET_B(_0279_),
    .Q(\second_row[5][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5503_ (.CLK(clknet_leaf_38_CLK),
    .D(_0814_),
    .RESET_B(_0280_),
    .Q(\second_row[5][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5504_ (.CLK(clknet_leaf_47_CLK),
    .D(_0815_),
    .RESET_B(_0281_),
    .Q(\second_row[5][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5505_ (.CLK(clknet_leaf_47_CLK),
    .D(_0816_),
    .RESET_B(_0282_),
    .Q(\second_row[5][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5506_ (.CLK(clknet_leaf_48_CLK),
    .D(_0817_),
    .RESET_B(_0283_),
    .Q(\second_row[5][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5507_ (.CLK(clknet_leaf_48_CLK),
    .D(_0818_),
    .RESET_B(_0284_),
    .Q(\second_row[5][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5508_ (.CLK(clknet_leaf_35_CLK),
    .D(_0819_),
    .RESET_B(_0285_),
    .Q(\second_row[6][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5509_ (.CLK(clknet_leaf_35_CLK),
    .D(_0820_),
    .RESET_B(_0286_),
    .Q(\second_row[6][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5510_ (.CLK(clknet_leaf_35_CLK),
    .D(_0821_),
    .RESET_B(_0287_),
    .Q(\second_row[6][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5511_ (.CLK(clknet_leaf_36_CLK),
    .D(_0822_),
    .RESET_B(_0288_),
    .Q(\second_row[6][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5512_ (.CLK(clknet_leaf_44_CLK),
    .D(_0823_),
    .RESET_B(_0289_),
    .Q(\second_row[6][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5513_ (.CLK(clknet_leaf_47_CLK),
    .D(_0824_),
    .RESET_B(_0290_),
    .Q(\second_row[6][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5514_ (.CLK(clknet_leaf_44_CLK),
    .D(_0825_),
    .RESET_B(_0291_),
    .Q(\second_row[6][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5515_ (.CLK(clknet_leaf_44_CLK),
    .D(_0826_),
    .RESET_B(_0292_),
    .Q(\second_row[6][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5516_ (.CLK(clknet_leaf_30_CLK),
    .D(_0827_),
    .RESET_B(_0293_),
    .Q(\second_row[7][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5517_ (.CLK(clknet_leaf_30_CLK),
    .D(_0828_),
    .RESET_B(_0294_),
    .Q(\second_row[7][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5518_ (.CLK(clknet_leaf_24_CLK),
    .D(_0829_),
    .RESET_B(_0295_),
    .Q(\second_row[7][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5519_ (.CLK(clknet_leaf_22_CLK),
    .D(_0830_),
    .RESET_B(_0296_),
    .Q(\second_row[7][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5520_ (.CLK(clknet_leaf_21_CLK),
    .D(_0831_),
    .RESET_B(_0297_),
    .Q(\second_row[7][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5521_ (.CLK(clknet_leaf_8_CLK),
    .D(_0832_),
    .RESET_B(_0298_),
    .Q(\second_row[7][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5522_ (.CLK(clknet_leaf_7_CLK),
    .D(_0833_),
    .RESET_B(_0299_),
    .Q(\second_row[7][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5523_ (.CLK(clknet_leaf_6_CLK),
    .D(_0834_),
    .RESET_B(_0300_),
    .Q(\second_row[7][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5524_ (.CLK(clknet_leaf_23_CLK),
    .D(_0835_),
    .RESET_B(_0301_),
    .Q(\second_row[8][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5525_ (.CLK(clknet_leaf_23_CLK),
    .D(_0836_),
    .RESET_B(_0302_),
    .Q(\second_row[8][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5526_ (.CLK(clknet_leaf_25_CLK),
    .D(_0837_),
    .RESET_B(_0303_),
    .Q(\second_row[8][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5527_ (.CLK(clknet_leaf_8_CLK),
    .D(_0838_),
    .RESET_B(_0304_),
    .Q(\second_row[8][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5528_ (.CLK(clknet_leaf_1_CLK),
    .D(_0839_),
    .RESET_B(_0305_),
    .Q(\second_row[8][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5529_ (.CLK(clknet_leaf_59_CLK),
    .D(_0840_),
    .RESET_B(_0306_),
    .Q(\second_row[8][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5530_ (.CLK(clknet_leaf_63_CLK),
    .D(_0841_),
    .RESET_B(_0307_),
    .Q(\second_row[8][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5531_ (.CLK(clknet_leaf_62_CLK),
    .D(_0842_),
    .RESET_B(_0308_),
    .Q(\second_row[8][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5532_ (.CLK(clknet_leaf_14_CLK),
    .D(_0843_),
    .RESET_B(_0309_),
    .Q(\second_row[9][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5533_ (.CLK(clknet_leaf_20_CLK),
    .D(_0844_),
    .RESET_B(_0310_),
    .Q(\second_row[9][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5534_ (.CLK(clknet_leaf_24_CLK),
    .D(_0845_),
    .RESET_B(_0311_),
    .Q(\second_row[9][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5535_ (.CLK(clknet_leaf_7_CLK),
    .D(_0846_),
    .RESET_B(_0312_),
    .Q(\second_row[9][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5536_ (.CLK(clknet_leaf_59_CLK),
    .D(_0847_),
    .RESET_B(_0313_),
    .Q(\second_row[9][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5537_ (.CLK(clknet_leaf_63_CLK),
    .D(_0848_),
    .RESET_B(_0314_),
    .Q(\second_row[9][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5538_ (.CLK(clknet_leaf_62_CLK),
    .D(_0849_),
    .RESET_B(_0315_),
    .Q(\second_row[9][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5539_ (.CLK(clknet_leaf_62_CLK),
    .D(_0850_),
    .RESET_B(_0316_),
    .Q(\second_row[9][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5540_ (.CLK(clknet_leaf_13_CLK),
    .D(_0851_),
    .RESET_B(_0317_),
    .Q(\second_row[10][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5541_ (.CLK(clknet_leaf_20_CLK),
    .D(_0852_),
    .RESET_B(_0318_),
    .Q(\second_row[10][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5542_ (.CLK(clknet_leaf_12_CLK),
    .D(_0853_),
    .RESET_B(_0319_),
    .Q(\second_row[10][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5543_ (.CLK(clknet_leaf_10_CLK),
    .D(_0854_),
    .RESET_B(_0320_),
    .Q(\second_row[10][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5544_ (.CLK(clknet_leaf_59_CLK),
    .D(_0855_),
    .RESET_B(_0321_),
    .Q(\second_row[10][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5545_ (.CLK(clknet_leaf_62_CLK),
    .D(_0856_),
    .RESET_B(_0322_),
    .Q(\second_row[10][5] ));
 sky130_fd_sc_hd__dfrtp_2 _5546_ (.CLK(clknet_leaf_62_CLK),
    .D(_0857_),
    .RESET_B(_0323_),
    .Q(\second_row[10][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5547_ (.CLK(clknet_leaf_62_CLK),
    .D(_0858_),
    .RESET_B(_0324_),
    .Q(\second_row[10][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5548_ (.CLK(clknet_leaf_15_CLK),
    .D(_0859_),
    .RESET_B(_0325_),
    .Q(\second_row[11][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5549_ (.CLK(clknet_leaf_16_CLK),
    .D(_0860_),
    .RESET_B(_0326_),
    .Q(\second_row[11][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5550_ (.CLK(clknet_leaf_12_CLK),
    .D(_0861_),
    .RESET_B(_0327_),
    .Q(\second_row[11][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5551_ (.CLK(clknet_leaf_11_CLK),
    .D(_0862_),
    .RESET_B(_0328_),
    .Q(\second_row[11][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5552_ (.CLK(clknet_leaf_2_CLK),
    .D(_0863_),
    .RESET_B(_0329_),
    .Q(\second_row[11][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5553_ (.CLK(clknet_leaf_11_CLK),
    .D(_0864_),
    .RESET_B(_0330_),
    .Q(\second_row[11][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5554_ (.CLK(clknet_leaf_3_CLK),
    .D(_0865_),
    .RESET_B(_0331_),
    .Q(\second_row[11][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5555_ (.CLK(clknet_leaf_2_CLK),
    .D(_0866_),
    .RESET_B(_0332_),
    .Q(\second_row[11][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5556_ (.CLK(clknet_leaf_16_CLK),
    .D(_0867_),
    .RESET_B(_0333_),
    .Q(\second_row[12][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5557_ (.CLK(clknet_leaf_16_CLK),
    .D(_0868_),
    .RESET_B(_0334_),
    .Q(\second_row[12][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5558_ (.CLK(clknet_leaf_15_CLK),
    .D(_0869_),
    .RESET_B(_0335_),
    .Q(\second_row[12][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5559_ (.CLK(clknet_leaf_9_CLK),
    .D(_0870_),
    .RESET_B(_0336_),
    .Q(\second_row[12][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5560_ (.CLK(clknet_leaf_5_CLK),
    .D(_0871_),
    .RESET_B(_0337_),
    .Q(\second_row[12][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5561_ (.CLK(clknet_leaf_63_CLK),
    .D(_0872_),
    .RESET_B(_0338_),
    .Q(\second_row[12][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5562_ (.CLK(clknet_leaf_63_CLK),
    .D(_0873_),
    .RESET_B(_0339_),
    .Q(\second_row[12][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5563_ (.CLK(clknet_leaf_63_CLK),
    .D(_0874_),
    .RESET_B(_0340_),
    .Q(\second_row[12][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5564_ (.CLK(clknet_leaf_23_CLK),
    .D(_0875_),
    .RESET_B(_0341_),
    .Q(\second_row[13][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5565_ (.CLK(clknet_leaf_23_CLK),
    .D(_0876_),
    .RESET_B(_0342_),
    .Q(\second_row[13][1] ));
 sky130_fd_sc_hd__dfrtp_2 _5566_ (.CLK(clknet_leaf_25_CLK),
    .D(_0877_),
    .RESET_B(_0343_),
    .Q(\second_row[13][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5567_ (.CLK(clknet_leaf_7_CLK),
    .D(_0878_),
    .RESET_B(_0344_),
    .Q(\second_row[13][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5568_ (.CLK(clknet_leaf_58_CLK),
    .D(_0879_),
    .RESET_B(_0345_),
    .Q(\second_row[13][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5569_ (.CLK(clknet_leaf_54_CLK),
    .D(_0880_),
    .RESET_B(_0346_),
    .Q(\second_row[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5570_ (.CLK(clknet_leaf_54_CLK),
    .D(_0881_),
    .RESET_B(_0347_),
    .Q(\second_row[13][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5571_ (.CLK(clknet_leaf_59_CLK),
    .D(_0882_),
    .RESET_B(_0348_),
    .Q(\second_row[13][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5572_ (.CLK(clknet_leaf_28_CLK),
    .D(_0883_),
    .RESET_B(_0349_),
    .Q(\second_row[14][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5573_ (.CLK(clknet_leaf_28_CLK),
    .D(_0884_),
    .RESET_B(_0350_),
    .Q(\second_row[14][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5574_ (.CLK(clknet_leaf_23_CLK),
    .D(_0885_),
    .RESET_B(_0351_),
    .Q(\second_row[14][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5575_ (.CLK(clknet_leaf_25_CLK),
    .D(_0886_),
    .RESET_B(_0352_),
    .Q(\second_row[14][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5576_ (.CLK(clknet_leaf_58_CLK),
    .D(_0887_),
    .RESET_B(_0353_),
    .Q(\second_row[14][4] ));
 sky130_fd_sc_hd__dfrtp_2 _5577_ (.CLK(clknet_leaf_59_CLK),
    .D(_0888_),
    .RESET_B(_0354_),
    .Q(\second_row[14][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5578_ (.CLK(clknet_leaf_62_CLK),
    .D(_0889_),
    .RESET_B(_0355_),
    .Q(\second_row[14][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5579_ (.CLK(clknet_leaf_62_CLK),
    .D(_0890_),
    .RESET_B(_0356_),
    .Q(\second_row[14][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5580_ (.CLK(clknet_leaf_28_CLK),
    .D(_0891_),
    .RESET_B(_0357_),
    .Q(\second_row[15][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5581_ (.CLK(clknet_leaf_23_CLK),
    .D(_0892_),
    .RESET_B(_0358_),
    .Q(\second_row[15][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5582_ (.CLK(clknet_leaf_24_CLK),
    .D(_0893_),
    .RESET_B(_0359_),
    .Q(\second_row[15][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5583_ (.CLK(clknet_leaf_7_CLK),
    .D(_0894_),
    .RESET_B(_0360_),
    .Q(\second_row[15][3] ));
 sky130_fd_sc_hd__dfrtp_2 _5584_ (.CLK(clknet_leaf_4_CLK),
    .D(_0895_),
    .RESET_B(_0361_),
    .Q(\second_row[15][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5585_ (.CLK(clknet_leaf_11_CLK),
    .D(_0896_),
    .RESET_B(_0362_),
    .Q(\second_row[15][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5586_ (.CLK(clknet_leaf_3_CLK),
    .D(_0897_),
    .RESET_B(_0363_),
    .Q(\second_row[15][6] ));
 sky130_fd_sc_hd__dfrtp_4 _5587_ (.CLK(clknet_leaf_1_CLK),
    .D(_0898_),
    .RESET_B(_0364_),
    .Q(\second_row[15][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5588_ (.CLK(clknet_leaf_14_CLK),
    .D(_0899_),
    .RESET_B(_0365_),
    .Q(\second_row[16][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5589_ (.CLK(clknet_leaf_14_CLK),
    .D(_0900_),
    .RESET_B(_0366_),
    .Q(\second_row[16][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5590_ (.CLK(clknet_leaf_12_CLK),
    .D(_0901_),
    .RESET_B(_0367_),
    .Q(\second_row[16][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5591_ (.CLK(clknet_leaf_11_CLK),
    .D(_0902_),
    .RESET_B(_0368_),
    .Q(\second_row[16][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5592_ (.CLK(clknet_leaf_2_CLK),
    .D(_0903_),
    .RESET_B(_0369_),
    .Q(\second_row[16][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5593_ (.CLK(clknet_leaf_11_CLK),
    .D(_0904_),
    .RESET_B(_0370_),
    .Q(\second_row[16][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5594_ (.CLK(clknet_leaf_5_CLK),
    .D(_0905_),
    .RESET_B(_0371_),
    .Q(\second_row[16][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5595_ (.CLK(clknet_leaf_5_CLK),
    .D(_0906_),
    .RESET_B(_0372_),
    .Q(\second_row[16][7] ));
 sky130_fd_sc_hd__dfrtp_4 _5596_ (.CLK(clknet_leaf_20_CLK),
    .D(_0907_),
    .RESET_B(_0373_),
    .Q(\second_row[17][0] ));
 sky130_fd_sc_hd__dfrtp_4 _5597_ (.CLK(clknet_leaf_20_CLK),
    .D(_0908_),
    .RESET_B(_0374_),
    .Q(\second_row[17][1] ));
 sky130_fd_sc_hd__dfrtp_4 _5598_ (.CLK(clknet_leaf_8_CLK),
    .D(_0909_),
    .RESET_B(_0375_),
    .Q(\second_row[17][2] ));
 sky130_fd_sc_hd__dfrtp_4 _5599_ (.CLK(clknet_leaf_10_CLK),
    .D(_0910_),
    .RESET_B(_0376_),
    .Q(\second_row[17][3] ));
 sky130_fd_sc_hd__dfrtp_4 _5600_ (.CLK(clknet_leaf_1_CLK),
    .D(_0911_),
    .RESET_B(_0377_),
    .Q(\second_row[17][4] ));
 sky130_fd_sc_hd__dfrtp_4 _5601_ (.CLK(clknet_leaf_4_CLK),
    .D(_0912_),
    .RESET_B(_0378_),
    .Q(\second_row[17][5] ));
 sky130_fd_sc_hd__dfrtp_4 _5602_ (.CLK(clknet_leaf_5_CLK),
    .D(_0913_),
    .RESET_B(_0379_),
    .Q(\second_row[17][6] ));
 sky130_fd_sc_hd__dfrtp_2 _5603_ (.CLK(clknet_leaf_5_CLK),
    .D(_0914_),
    .RESET_B(_0380_),
    .Q(\second_row[17][7] ));
 sky130_fd_sc_hd__dfrtp_2 _5604_ (.CLK(clknet_leaf_12_CLK),
    .D(_0915_),
    .RESET_B(_0381_),
    .Q(\third_row[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5605_ (.CLK(clknet_leaf_8_CLK),
    .D(_0916_),
    .RESET_B(_0382_),
    .Q(\third_row[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5606_ (.CLK(clknet_leaf_12_CLK),
    .D(_0917_),
    .RESET_B(_0383_),
    .Q(\third_row[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5607_ (.CLK(clknet_leaf_3_CLK),
    .D(_0918_),
    .RESET_B(_0384_),
    .Q(\third_row[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5608_ (.CLK(clknet_leaf_2_CLK),
    .D(_0919_),
    .RESET_B(_0385_),
    .Q(\third_row[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5609_ (.CLK(clknet_leaf_64_CLK),
    .D(_0920_),
    .RESET_B(_0386_),
    .Q(\third_row[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5610_ (.CLK(clknet_leaf_51_CLK),
    .D(_0921_),
    .RESET_B(_0387_),
    .Q(\third_row[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5611_ (.CLK(clknet_leaf_64_CLK),
    .D(_0922_),
    .RESET_B(_0388_),
    .Q(\third_row[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5612_ (.CLK(clknet_leaf_41_CLK),
    .D(_0923_),
    .RESET_B(_0389_),
    .Q(\third_row[1][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5613_ (.CLK(clknet_leaf_36_CLK),
    .D(_0924_),
    .RESET_B(_0390_),
    .Q(\third_row[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5614_ (.CLK(clknet_leaf_43_CLK),
    .D(_0925_),
    .RESET_B(_0391_),
    .Q(\third_row[1][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5615_ (.CLK(clknet_leaf_43_CLK),
    .D(_0926_),
    .RESET_B(_0392_),
    .Q(\third_row[1][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5616_ (.CLK(clknet_leaf_57_CLK),
    .D(_0927_),
    .RESET_B(_0393_),
    .Q(\third_row[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5617_ (.CLK(clknet_leaf_51_CLK),
    .D(_0928_),
    .RESET_B(_0394_),
    .Q(\third_row[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5618_ (.CLK(clknet_leaf_52_CLK),
    .D(_0929_),
    .RESET_B(_0395_),
    .Q(\third_row[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5619_ (.CLK(clknet_leaf_60_CLK),
    .D(_0930_),
    .RESET_B(_0396_),
    .Q(\third_row[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5620_ (.CLK(clknet_leaf_41_CLK),
    .D(_0931_),
    .RESET_B(_0397_),
    .Q(\third_row[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5621_ (.CLK(clknet_leaf_41_CLK),
    .D(_0932_),
    .RESET_B(_0398_),
    .Q(\third_row[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5622_ (.CLK(clknet_leaf_26_CLK),
    .D(_0933_),
    .RESET_B(_0399_),
    .Q(\third_row[2][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5623_ (.CLK(clknet_leaf_45_CLK),
    .D(_0934_),
    .RESET_B(_0400_),
    .Q(\third_row[2][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5624_ (.CLK(clknet_leaf_56_CLK),
    .D(_0935_),
    .RESET_B(_0401_),
    .Q(\third_row[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5625_ (.CLK(clknet_leaf_55_CLK),
    .D(_0936_),
    .RESET_B(_0402_),
    .Q(\third_row[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5626_ (.CLK(clknet_leaf_54_CLK),
    .D(_0937_),
    .RESET_B(_0403_),
    .Q(\third_row[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5627_ (.CLK(clknet_leaf_60_CLK),
    .D(_0938_),
    .RESET_B(_0404_),
    .Q(\third_row[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5628_ (.CLK(clknet_leaf_41_CLK),
    .D(_0939_),
    .RESET_B(_0405_),
    .Q(\third_row[3][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5629_ (.CLK(clknet_leaf_39_CLK),
    .D(_0940_),
    .RESET_B(_0406_),
    .Q(\third_row[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5630_ (.CLK(clknet_leaf_26_CLK),
    .D(_0941_),
    .RESET_B(_0407_),
    .Q(\third_row[3][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5631_ (.CLK(clknet_leaf_42_CLK),
    .D(_0942_),
    .RESET_B(_0408_),
    .Q(\third_row[3][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5632_ (.CLK(clknet_leaf_56_CLK),
    .D(_0943_),
    .RESET_B(_0409_),
    .Q(\third_row[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5633_ (.CLK(clknet_leaf_50_CLK),
    .D(_0944_),
    .RESET_B(_0410_),
    .Q(\third_row[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5634_ (.CLK(clknet_leaf_49_CLK),
    .D(_0945_),
    .RESET_B(_0411_),
    .Q(\third_row[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5635_ (.CLK(clknet_leaf_60_CLK),
    .D(_0946_),
    .RESET_B(_0412_),
    .Q(\third_row[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5636_ (.CLK(clknet_leaf_42_CLK),
    .D(_0947_),
    .RESET_B(_0413_),
    .Q(\third_row[4][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5637_ (.CLK(clknet_leaf_39_CLK),
    .D(_0948_),
    .RESET_B(_0414_),
    .Q(\third_row[4][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5638_ (.CLK(clknet_leaf_42_CLK),
    .D(_0949_),
    .RESET_B(_0415_),
    .Q(\third_row[4][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5639_ (.CLK(clknet_leaf_45_CLK),
    .D(_0950_),
    .RESET_B(_0416_),
    .Q(\third_row[4][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5640_ (.CLK(clknet_leaf_45_CLK),
    .D(_0951_),
    .RESET_B(_0417_),
    .Q(\third_row[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5641_ (.CLK(clknet_leaf_49_CLK),
    .D(_0952_),
    .RESET_B(_0418_),
    .Q(\third_row[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5642_ (.CLK(clknet_leaf_49_CLK),
    .D(_0953_),
    .RESET_B(_0419_),
    .Q(\third_row[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5643_ (.CLK(clknet_leaf_49_CLK),
    .D(_0954_),
    .RESET_B(_0420_),
    .Q(\third_row[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5644_ (.CLK(clknet_leaf_39_CLK),
    .D(_0955_),
    .RESET_B(_0421_),
    .Q(\third_row[5][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5645_ (.CLK(clknet_leaf_39_CLK),
    .D(_0956_),
    .RESET_B(_0422_),
    .Q(\third_row[5][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5646_ (.CLK(clknet_leaf_45_CLK),
    .D(_0957_),
    .RESET_B(_0423_),
    .Q(\third_row[5][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5647_ (.CLK(clknet_leaf_45_CLK),
    .D(_0958_),
    .RESET_B(_0424_),
    .Q(\third_row[5][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5648_ (.CLK(clknet_leaf_46_CLK),
    .D(_0959_),
    .RESET_B(_0425_),
    .Q(\third_row[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5649_ (.CLK(clknet_leaf_47_CLK),
    .D(_0960_),
    .RESET_B(_0426_),
    .Q(\third_row[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5650_ (.CLK(clknet_leaf_49_CLK),
    .D(_0961_),
    .RESET_B(_0427_),
    .Q(\third_row[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5651_ (.CLK(clknet_leaf_48_CLK),
    .D(_0962_),
    .RESET_B(_0428_),
    .Q(\third_row[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5652_ (.CLK(clknet_leaf_39_CLK),
    .D(_0963_),
    .RESET_B(_0429_),
    .Q(\third_row[6][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5653_ (.CLK(clknet_leaf_39_CLK),
    .D(_0964_),
    .RESET_B(_0430_),
    .Q(\third_row[6][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5654_ (.CLK(clknet_leaf_46_CLK),
    .D(_0965_),
    .RESET_B(_0431_),
    .Q(\third_row[6][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5655_ (.CLK(clknet_leaf_45_CLK),
    .D(_0966_),
    .RESET_B(_0432_),
    .Q(\third_row[6][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5656_ (.CLK(clknet_leaf_46_CLK),
    .D(_0967_),
    .RESET_B(_0433_),
    .Q(\third_row[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5657_ (.CLK(clknet_leaf_47_CLK),
    .D(_0968_),
    .RESET_B(_0434_),
    .Q(\third_row[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5658_ (.CLK(clknet_leaf_49_CLK),
    .D(_0969_),
    .RESET_B(_0435_),
    .Q(\third_row[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5659_ (.CLK(clknet_leaf_49_CLK),
    .D(_0970_),
    .RESET_B(_0436_),
    .Q(\third_row[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5660_ (.CLK(clknet_leaf_41_CLK),
    .D(_0971_),
    .RESET_B(_0437_),
    .Q(\third_row[7][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5661_ (.CLK(clknet_leaf_40_CLK),
    .D(_0972_),
    .RESET_B(_0438_),
    .Q(\third_row[7][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5662_ (.CLK(clknet_leaf_45_CLK),
    .D(_0973_),
    .RESET_B(_0439_),
    .Q(\third_row[7][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5663_ (.CLK(clknet_leaf_43_CLK),
    .D(_0974_),
    .RESET_B(_0440_),
    .Q(\third_row[7][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5664_ (.CLK(clknet_leaf_56_CLK),
    .D(_0975_),
    .RESET_B(_0441_),
    .Q(\third_row[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5665_ (.CLK(clknet_leaf_54_CLK),
    .D(_0976_),
    .RESET_B(_0442_),
    .Q(\third_row[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5666_ (.CLK(clknet_leaf_52_CLK),
    .D(_0977_),
    .RESET_B(_0443_),
    .Q(\third_row[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5667_ (.CLK(clknet_leaf_60_CLK),
    .D(_0978_),
    .RESET_B(_0444_),
    .Q(\third_row[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5668_ (.CLK(clknet_leaf_41_CLK),
    .D(_0979_),
    .RESET_B(_0445_),
    .Q(\third_row[8][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5669_ (.CLK(clknet_leaf_41_CLK),
    .D(_0980_),
    .RESET_B(_0446_),
    .Q(\third_row[8][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5670_ (.CLK(clknet_leaf_26_CLK),
    .D(_0981_),
    .RESET_B(_0447_),
    .Q(\third_row[8][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5671_ (.CLK(clknet_leaf_61_CLK),
    .D(_0982_),
    .RESET_B(_0448_),
    .Q(\third_row[8][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5672_ (.CLK(clknet_leaf_56_CLK),
    .D(_0983_),
    .RESET_B(_0449_),
    .Q(\third_row[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5673_ (.CLK(clknet_leaf_55_CLK),
    .D(_0984_),
    .RESET_B(_0450_),
    .Q(\third_row[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5674_ (.CLK(clknet_leaf_53_CLK),
    .D(_0985_),
    .RESET_B(_0451_),
    .Q(\third_row[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5675_ (.CLK(clknet_leaf_53_CLK),
    .D(_0986_),
    .RESET_B(_0452_),
    .Q(\third_row[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5676_ (.CLK(clknet_leaf_42_CLK),
    .D(_0987_),
    .RESET_B(_0453_),
    .Q(\third_row[9][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5677_ (.CLK(clknet_leaf_39_CLK),
    .D(_0988_),
    .RESET_B(_0454_),
    .Q(\third_row[9][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5678_ (.CLK(clknet_leaf_42_CLK),
    .D(_0989_),
    .RESET_B(_0455_),
    .Q(\third_row[9][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5679_ (.CLK(clknet_leaf_51_CLK),
    .D(_0990_),
    .RESET_B(_0456_),
    .Q(\third_row[9][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5680_ (.CLK(clknet_leaf_56_CLK),
    .D(_0991_),
    .RESET_B(_0457_),
    .Q(\third_row[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5681_ (.CLK(clknet_leaf_49_CLK),
    .D(_0992_),
    .RESET_B(_0458_),
    .Q(\third_row[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5682_ (.CLK(clknet_leaf_49_CLK),
    .D(_0993_),
    .RESET_B(_0459_),
    .Q(\third_row[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5683_ (.CLK(clknet_leaf_53_CLK),
    .D(_0994_),
    .RESET_B(_0460_),
    .Q(\third_row[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5684_ (.CLK(clknet_leaf_39_CLK),
    .D(_0995_),
    .RESET_B(_0461_),
    .Q(\third_row[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5685_ (.CLK(clknet_leaf_39_CLK),
    .D(_0996_),
    .RESET_B(_0462_),
    .Q(\third_row[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5686_ (.CLK(clknet_leaf_26_CLK),
    .D(_0997_),
    .RESET_B(_0463_),
    .Q(\third_row[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5687_ (.CLK(clknet_leaf_56_CLK),
    .D(_0998_),
    .RESET_B(_0464_),
    .Q(\third_row[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5688_ (.CLK(clknet_leaf_56_CLK),
    .D(_0999_),
    .RESET_B(_0465_),
    .Q(\third_row[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5689_ (.CLK(clknet_leaf_54_CLK),
    .D(_1000_),
    .RESET_B(_0466_),
    .Q(\third_row[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5690_ (.CLK(clknet_leaf_53_CLK),
    .D(_1001_),
    .RESET_B(_0467_),
    .Q(\third_row[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5691_ (.CLK(clknet_leaf_53_CLK),
    .D(_1002_),
    .RESET_B(_0468_),
    .Q(\third_row[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5692_ (.CLK(clknet_leaf_40_CLK),
    .D(_1003_),
    .RESET_B(_0469_),
    .Q(\third_row[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5693_ (.CLK(clknet_leaf_40_CLK),
    .D(_1004_),
    .RESET_B(_0470_),
    .Q(\third_row[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5694_ (.CLK(clknet_leaf_26_CLK),
    .D(_1005_),
    .RESET_B(_0471_),
    .Q(\third_row[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5695_ (.CLK(clknet_leaf_58_CLK),
    .D(_1006_),
    .RESET_B(_0472_),
    .Q(\third_row[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5696_ (.CLK(clknet_leaf_56_CLK),
    .D(_1007_),
    .RESET_B(_0473_),
    .Q(\third_row[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5697_ (.CLK(clknet_leaf_49_CLK),
    .D(_1008_),
    .RESET_B(_0474_),
    .Q(\third_row[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5698_ (.CLK(clknet_leaf_52_CLK),
    .D(_1009_),
    .RESET_B(_0475_),
    .Q(\third_row[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5699_ (.CLK(clknet_leaf_60_CLK),
    .D(_1010_),
    .RESET_B(_0476_),
    .Q(\third_row[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5700_ (.CLK(clknet_leaf_41_CLK),
    .D(_1011_),
    .RESET_B(_0477_),
    .Q(\third_row[12][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5701_ (.CLK(clknet_leaf_39_CLK),
    .D(_1012_),
    .RESET_B(_0478_),
    .Q(\third_row[12][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5702_ (.CLK(clknet_leaf_42_CLK),
    .D(_1013_),
    .RESET_B(_0479_),
    .Q(\third_row[12][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5703_ (.CLK(clknet_leaf_53_CLK),
    .D(_1014_),
    .RESET_B(_0480_),
    .Q(\third_row[12][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5704_ (.CLK(clknet_leaf_56_CLK),
    .D(_1015_),
    .RESET_B(_0481_),
    .Q(\third_row[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5705_ (.CLK(clknet_leaf_49_CLK),
    .D(_1016_),
    .RESET_B(_0482_),
    .Q(\third_row[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5706_ (.CLK(clknet_leaf_53_CLK),
    .D(_1017_),
    .RESET_B(_0483_),
    .Q(\third_row[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5707_ (.CLK(clknet_leaf_53_CLK),
    .D(_1018_),
    .RESET_B(_0484_),
    .Q(\third_row[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5708_ (.CLK(clknet_leaf_39_CLK),
    .D(_1019_),
    .RESET_B(_0485_),
    .Q(\third_row[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5709_ (.CLK(clknet_leaf_45_CLK),
    .D(_1020_),
    .RESET_B(_0486_),
    .Q(\third_row[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5710_ (.CLK(clknet_leaf_42_CLK),
    .D(_1021_),
    .RESET_B(_0487_),
    .Q(\third_row[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5711_ (.CLK(clknet_leaf_61_CLK),
    .D(_1022_),
    .RESET_B(_0488_),
    .Q(\third_row[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5712_ (.CLK(clknet_leaf_43_CLK),
    .D(_1023_),
    .RESET_B(_0489_),
    .Q(\third_row[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5713_ (.CLK(clknet_leaf_49_CLK),
    .D(_1024_),
    .RESET_B(_0490_),
    .Q(\third_row[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5714_ (.CLK(clknet_leaf_53_CLK),
    .D(_1025_),
    .RESET_B(_0491_),
    .Q(\third_row[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5715_ (.CLK(clknet_leaf_53_CLK),
    .D(_1026_),
    .RESET_B(_0492_),
    .Q(\third_row[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5716_ (.CLK(clknet_leaf_43_CLK),
    .D(_1027_),
    .RESET_B(_0493_),
    .Q(\third_row[14][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5717_ (.CLK(clknet_leaf_43_CLK),
    .D(_1028_),
    .RESET_B(_0494_),
    .Q(\third_row[14][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5718_ (.CLK(clknet_leaf_43_CLK),
    .D(_1029_),
    .RESET_B(_0495_),
    .Q(\third_row[14][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5719_ (.CLK(clknet_leaf_43_CLK),
    .D(_1030_),
    .RESET_B(_0496_),
    .Q(\third_row[14][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5720_ (.CLK(clknet_leaf_44_CLK),
    .D(_1031_),
    .RESET_B(_0497_),
    .Q(\third_row[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5721_ (.CLK(clknet_leaf_50_CLK),
    .D(_1032_),
    .RESET_B(_0498_),
    .Q(\third_row[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5722_ (.CLK(clknet_leaf_51_CLK),
    .D(_1033_),
    .RESET_B(_0499_),
    .Q(\third_row[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5723_ (.CLK(clknet_leaf_53_CLK),
    .D(_1034_),
    .RESET_B(_0500_),
    .Q(\third_row[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5724_ (.CLK(clknet_leaf_40_CLK),
    .D(_1035_),
    .RESET_B(_0501_),
    .Q(\third_row[15][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5725_ (.CLK(clknet_leaf_40_CLK),
    .D(_1036_),
    .RESET_B(_0502_),
    .Q(\third_row[15][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5726_ (.CLK(clknet_leaf_42_CLK),
    .D(_1037_),
    .RESET_B(_0503_),
    .Q(\third_row[15][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5727_ (.CLK(clknet_leaf_43_CLK),
    .D(_1038_),
    .RESET_B(_0504_),
    .Q(\third_row[15][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5728_ (.CLK(clknet_leaf_57_CLK),
    .D(_1039_),
    .RESET_B(_0505_),
    .Q(\third_row[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5729_ (.CLK(clknet_leaf_55_CLK),
    .D(_1040_),
    .RESET_B(_0506_),
    .Q(\third_row[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5730_ (.CLK(clknet_leaf_52_CLK),
    .D(_1041_),
    .RESET_B(_0507_),
    .Q(\third_row[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5731_ (.CLK(clknet_leaf_61_CLK),
    .D(_1042_),
    .RESET_B(_0508_),
    .Q(\third_row[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5732_ (.CLK(clknet_3_6__leaf_CLK),
    .D(_1043_),
    .RESET_B(_0509_),
    .Q(\third_row[16][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5733_ (.CLK(clknet_leaf_41_CLK),
    .D(_1044_),
    .RESET_B(_0510_),
    .Q(\third_row[16][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5734_ (.CLK(clknet_leaf_25_CLK),
    .D(_1045_),
    .RESET_B(_0511_),
    .Q(\third_row[16][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5735_ (.CLK(clknet_leaf_57_CLK),
    .D(_1046_),
    .RESET_B(_0512_),
    .Q(\third_row[16][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5736_ (.CLK(clknet_leaf_56_CLK),
    .D(_1047_),
    .RESET_B(_0513_),
    .Q(\third_row[16][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5737_ (.CLK(clknet_leaf_52_CLK),
    .D(_1048_),
    .RESET_B(_0514_),
    .Q(\third_row[16][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5738_ (.CLK(clknet_leaf_50_CLK),
    .D(_1049_),
    .RESET_B(_0515_),
    .Q(\third_row[16][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5739_ (.CLK(clknet_leaf_60_CLK),
    .D(_1050_),
    .RESET_B(_0516_),
    .Q(\third_row[16][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5740_ (.CLK(clknet_leaf_15_CLK),
    .D(_1051_),
    .RESET_B(_0517_),
    .Q(\first_row[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5741_ (.CLK(clknet_leaf_15_CLK),
    .D(_1052_),
    .RESET_B(_0518_),
    .Q(\first_row[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5742_ (.CLK(clknet_leaf_12_CLK),
    .D(_1053_),
    .RESET_B(_0519_),
    .Q(\first_row[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5743_ (.CLK(clknet_leaf_12_CLK),
    .D(_1054_),
    .RESET_B(_0520_),
    .Q(\first_row[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5744_ (.CLK(clknet_leaf_2_CLK),
    .D(_1055_),
    .RESET_B(_0521_),
    .Q(\first_row[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5745_ (.CLK(clknet_leaf_64_CLK),
    .D(_1056_),
    .RESET_B(_0522_),
    .Q(\first_row[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5746_ (.CLK(clknet_leaf_64_CLK),
    .D(_1057_),
    .RESET_B(_0523_),
    .Q(\first_row[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5747_ (.CLK(clknet_leaf_64_CLK),
    .D(_1058_),
    .RESET_B(_0524_),
    .Q(\first_row[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5748_ (.CLK(clknet_leaf_42_CLK),
    .D(_1059_),
    .RESET_B(_0525_),
    .Q(\third_row[17][0] ));
 sky130_fd_sc_hd__dfrtp_1 _5749_ (.CLK(clknet_leaf_41_CLK),
    .D(_1060_),
    .RESET_B(_0526_),
    .Q(\third_row[17][1] ));
 sky130_fd_sc_hd__dfrtp_1 _5750_ (.CLK(clknet_leaf_42_CLK),
    .D(_1061_),
    .RESET_B(_0527_),
    .Q(\third_row[17][2] ));
 sky130_fd_sc_hd__dfrtp_1 _5751_ (.CLK(clknet_leaf_61_CLK),
    .D(_1062_),
    .RESET_B(_0528_),
    .Q(\third_row[17][3] ));
 sky130_fd_sc_hd__dfrtp_1 _5752_ (.CLK(clknet_leaf_53_CLK),
    .D(_1063_),
    .RESET_B(_0529_),
    .Q(\third_row[17][4] ));
 sky130_fd_sc_hd__dfrtp_1 _5753_ (.CLK(clknet_leaf_52_CLK),
    .D(_1064_),
    .RESET_B(_0530_),
    .Q(\third_row[17][5] ));
 sky130_fd_sc_hd__dfrtp_1 _5754_ (.CLK(clknet_leaf_50_CLK),
    .D(_1065_),
    .RESET_B(_0531_),
    .Q(\third_row[17][6] ));
 sky130_fd_sc_hd__dfrtp_1 _5755_ (.CLK(clknet_leaf_60_CLK),
    .D(_1066_),
    .RESET_B(_0532_),
    .Q(\third_row[17][7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1207 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(pixel_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(pixel_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(pixel_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(pixel_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(pixel_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(pixel_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(pixel_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_8 input8 (.A(pixel_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(rst),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(valid_in),
    .X(net10));
 sky130_fd_sc_hd__buf_1 output11 (.A(net11),
    .X(pixel_out[0]));
 sky130_fd_sc_hd__buf_1 output12 (.A(net12),
    .X(pixel_out[1]));
 sky130_fd_sc_hd__buf_1 output13 (.A(net13),
    .X(pixel_out[2]));
 sky130_fd_sc_hd__buf_1 output14 (.A(net14),
    .X(pixel_out[3]));
 sky130_fd_sc_hd__buf_1 output15 (.A(net15),
    .X(pixel_out[4]));
 sky130_fd_sc_hd__buf_1 output16 (.A(net16),
    .X(pixel_out[5]));
 sky130_fd_sc_hd__buf_1 output17 (.A(net17),
    .X(pixel_out[6]));
 sky130_fd_sc_hd__buf_1 output18 (.A(net18),
    .X(pixel_out[7]));
 sky130_fd_sc_hd__buf_1 output19 (.A(net19),
    .X(valid_out));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_6_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_7_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_16_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_CLK (.A(clknet_3_2__leaf_CLK),
    .X(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_CLK (.A(clknet_3_3__leaf_CLK),
    .X(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_38_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_CLK (.A(clknet_3_7__leaf_CLK),
    .X(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_CLK (.A(clknet_3_6__leaf_CLK),
    .X(clknet_leaf_41_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_CLK (.A(clknet_3_5__leaf_CLK),
    .X(clknet_leaf_49_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_53_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_CLK (.A(clknet_3_4__leaf_CLK),
    .X(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_CLK (.A(clknet_3_1__leaf_CLK),
    .X(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_62_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_CLK (.A(clknet_3_0__leaf_CLK),
    .X(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_1__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_2__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_3__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_4__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_5__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_6__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_CLK (.A(clknet_0_CLK),
    .X(clknet_3_7__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_3_0__leaf_CLK));
 sky130_fd_sc_hd__inv_12 clkload1 (.A(clknet_3_1__leaf_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_3_3__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_4__leaf_CLK));
 sky130_fd_sc_hd__inv_12 clkload4 (.A(clknet_3_5__leaf_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload5 (.A(clknet_3_6__leaf_CLK));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_7__leaf_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload7 (.A(clknet_leaf_0_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_1_CLK));
 sky130_fd_sc_hd__inv_6 clkload9 (.A(clknet_leaf_2_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_leaf_3_CLK));
 sky130_fd_sc_hd__clkinv_8 clkload11 (.A(clknet_leaf_4_CLK));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_leaf_5_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload13 (.A(clknet_leaf_63_CLK));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_leaf_64_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload15 (.A(clknet_leaf_57_CLK));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_58_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload17 (.A(clknet_leaf_59_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_60_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload19 (.A(clknet_leaf_61_CLK));
 sky130_fd_sc_hd__clkbuf_4 clkload20 (.A(clknet_leaf_8_CLK));
 sky130_fd_sc_hd__inv_6 clkload21 (.A(clknet_leaf_9_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload22 (.A(clknet_leaf_10_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload23 (.A(clknet_leaf_11_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload24 (.A(clknet_leaf_12_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload25 (.A(clknet_leaf_13_CLK));
 sky130_fd_sc_hd__inv_6 clkload26 (.A(clknet_leaf_14_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload27 (.A(clknet_leaf_15_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload28 (.A(clknet_leaf_17_CLK));
 sky130_fd_sc_hd__inv_6 clkload29 (.A(clknet_leaf_18_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload30 (.A(clknet_leaf_19_CLK));
 sky130_fd_sc_hd__clkbuf_4 clkload31 (.A(clknet_leaf_20_CLK));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_21_CLK));
 sky130_fd_sc_hd__clkbuf_4 clkload33 (.A(clknet_leaf_22_CLK));
 sky130_fd_sc_hd__clkinvlp_2 clkload34 (.A(clknet_leaf_23_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload35 (.A(clknet_leaf_24_CLK));
 sky130_fd_sc_hd__inv_6 clkload36 (.A(clknet_leaf_25_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload37 (.A(clknet_leaf_42_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload38 (.A(clknet_leaf_43_CLK));
 sky130_fd_sc_hd__inv_6 clkload39 (.A(clknet_leaf_50_CLK));
 sky130_fd_sc_hd__inv_6 clkload40 (.A(clknet_leaf_51_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload41 (.A(clknet_leaf_52_CLK));
 sky130_fd_sc_hd__inv_6 clkload42 (.A(clknet_leaf_54_CLK));
 sky130_fd_sc_hd__inv_6 clkload43 (.A(clknet_leaf_55_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload44 (.A(clknet_leaf_56_CLK));
 sky130_fd_sc_hd__clkinvlp_2 clkload45 (.A(clknet_leaf_44_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload46 (.A(clknet_leaf_45_CLK));
 sky130_fd_sc_hd__inv_8 clkload47 (.A(clknet_leaf_46_CLK));
 sky130_fd_sc_hd__clkbuf_4 clkload48 (.A(clknet_leaf_47_CLK));
 sky130_fd_sc_hd__inv_8 clkload49 (.A(clknet_leaf_48_CLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload50 (.A(clknet_leaf_26_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload51 (.A(clknet_leaf_28_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload52 (.A(clknet_leaf_29_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload53 (.A(clknet_leaf_30_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload54 (.A(clknet_leaf_40_CLK));
 sky130_fd_sc_hd__inv_8 clkload55 (.A(clknet_leaf_31_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload56 (.A(clknet_leaf_32_CLK));
 sky130_fd_sc_hd__clkinv_1 clkload57 (.A(clknet_leaf_33_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload58 (.A(clknet_leaf_34_CLK));
 sky130_fd_sc_hd__clkinv_4 clkload59 (.A(clknet_leaf_35_CLK));
 sky130_fd_sc_hd__inv_8 clkload60 (.A(clknet_leaf_36_CLK));
 sky130_fd_sc_hd__inv_6 clkload61 (.A(clknet_leaf_37_CLK));
 sky130_fd_sc_hd__bufinv_16 clkload62 (.A(clknet_leaf_39_CLK));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\second_row[10][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\second_row[15][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\second_row[15][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\second_row[16][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\second_row[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\second_row[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\second_row[9][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\second_row[9][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_2286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net5));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_583 ();
endmodule
